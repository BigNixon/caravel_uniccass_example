// This is the unpowered netlist.
module wb_buttons_leds (buttons,
    clk,
    i_wb_cyc,
    i_wb_stb,
    i_wb_we,
    o_wb_ack,
    o_wb_stall,
    reset,
    i_wb_addr,
    i_wb_data,
    led_enb,
    leds,
    o_wb_data);
 input buttons;
 input clk;
 input i_wb_cyc;
 input i_wb_stb;
 input i_wb_we;
 output o_wb_ack;
 output o_wb_stall;
 input reset;
 input [31:0] i_wb_addr;
 input [31:0] i_wb_data;
 output [11:0] led_enb;
 output [11:0] leds;
 output [31:0] o_wb_data;

 wire net939;
 wire net949;
 wire net950;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net951;
 wire \ApproximateM_inst.lob_16.lob1.genblk1[10].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob1.genblk1[11].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob1.genblk1[12].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob1.genblk1[13].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob1.genblk1[14].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob1.genblk1[1].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob1.genblk1[2].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob1.genblk1[3].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob1.genblk1[4].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob1.genblk1[5].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob1.genblk1[6].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob1.genblk1[7].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob1.genblk1[8].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob1.genblk1[9].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob1.genblk2.mux_final.sel ;
 wire \ApproximateM_inst.lob_16.lob1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob2.genblk1[10].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob2.genblk1[11].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob2.genblk1[12].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob2.genblk1[13].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob2.genblk1[14].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob2.genblk1[1].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob2.genblk1[2].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob2.genblk1[3].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob2.genblk1[4].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob2.genblk1[5].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob2.genblk1[6].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob2.genblk1[7].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob2.genblk1[8].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob2.genblk1[9].genblk1.mux.sel ;
 wire \ApproximateM_inst.lob_16.lob2.genblk2.mux_final.sel ;
 wire \ApproximateM_inst.lob_16.lob2.mux.sel ;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire \cla_inst.in1[16] ;
 wire \cla_inst.in1[17] ;
 wire \cla_inst.in1[18] ;
 wire \cla_inst.in1[19] ;
 wire \cla_inst.in1[20] ;
 wire \cla_inst.in1[21] ;
 wire \cla_inst.in1[22] ;
 wire \cla_inst.in1[23] ;
 wire \cla_inst.in1[24] ;
 wire \cla_inst.in1[25] ;
 wire \cla_inst.in1[26] ;
 wire \cla_inst.in1[27] ;
 wire \cla_inst.in1[28] ;
 wire \cla_inst.in1[29] ;
 wire \cla_inst.in1[30] ;
 wire \cla_inst.in1[31] ;
 wire \cla_inst.in2[16] ;
 wire \cla_inst.in2[17] ;
 wire \cla_inst.in2[18] ;
 wire \cla_inst.in2[19] ;
 wire \cla_inst.in2[20] ;
 wire \cla_inst.in2[21] ;
 wire \cla_inst.in2[22] ;
 wire \cla_inst.in2[23] ;
 wire \cla_inst.in2[24] ;
 wire \cla_inst.in2[25] ;
 wire \cla_inst.in2[26] ;
 wire \cla_inst.in2[27] ;
 wire \cla_inst.in2[28] ;
 wire \cla_inst.in2[29] ;
 wire \cla_inst.in2[30] ;
 wire \cla_inst.in2[31] ;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \op_code[0] ;
 wire \op_code[1] ;
 wire \op_code[2] ;
 wire \op_code[3] ;
 wire \salida[0] ;
 wire \salida[10] ;
 wire \salida[11] ;
 wire \salida[12] ;
 wire \salida[13] ;
 wire \salida[14] ;
 wire \salida[15] ;
 wire \salida[16] ;
 wire \salida[17] ;
 wire \salida[18] ;
 wire \salida[19] ;
 wire \salida[1] ;
 wire \salida[20] ;
 wire \salida[21] ;
 wire \salida[22] ;
 wire \salida[23] ;
 wire \salida[24] ;
 wire \salida[25] ;
 wire \salida[26] ;
 wire \salida[27] ;
 wire \salida[28] ;
 wire \salida[29] ;
 wire \salida[2] ;
 wire \salida[30] ;
 wire \salida[31] ;
 wire \salida[32] ;
 wire \salida[33] ;
 wire \salida[34] ;
 wire \salida[35] ;
 wire \salida[36] ;
 wire \salida[37] ;
 wire \salida[38] ;
 wire \salida[39] ;
 wire \salida[3] ;
 wire \salida[40] ;
 wire \salida[41] ;
 wire \salida[42] ;
 wire \salida[43] ;
 wire \salida[44] ;
 wire \salida[45] ;
 wire \salida[46] ;
 wire \salida[47] ;
 wire \salida[48] ;
 wire \salida[49] ;
 wire \salida[4] ;
 wire \salida[50] ;
 wire \salida[51] ;
 wire \salida[52] ;
 wire \salida[53] ;
 wire \salida[54] ;
 wire \salida[55] ;
 wire \salida[56] ;
 wire \salida[57] ;
 wire \salida[58] ;
 wire \salida[59] ;
 wire \salida[5] ;
 wire \salida[60] ;
 wire \salida[61] ;
 wire \salida[62] ;
 wire \salida[63] ;
 wire \salida[6] ;
 wire \salida[7] ;
 wire \salida[8] ;
 wire \salida[9] ;
 wire \sel_op[0] ;
 wire \sel_op[1] ;
 wire \sel_op[2] ;
 wire \sel_op[3] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\ApproximateM_inst.lob_16.lob1.genblk1[9].genblk1.mux.sel ));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_05981_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_06732_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_08223_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_08692_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_08693_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(\cla_inst.in2[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_00100_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_00100_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_00100_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(_06047_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_00100_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(_06368_));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(_07624_));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(_07627_));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(\cla_inst.in1[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(\salida[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_00653_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_03527_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_03847_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_04764_));
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_842 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_926 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_899 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1066 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_930 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1064 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1064 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1098 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1068 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1064 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1048 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_871 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1016 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1039 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1059 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_960 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_644 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_972 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_984 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_703 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_898 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_980 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1003 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_927 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_868 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_989 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_4 _08717_ (.A(\ApproximateM_inst.lob_16.lob2.genblk1[7].genblk1.mux.sel ),
    .Y(_03182_));
 sky130_fd_sc_hd__clkinv_4 _08718_ (.A(net540),
    .Y(_03193_));
 sky130_fd_sc_hd__inv_2 _08719_ (.A(net559),
    .Y(_03203_));
 sky130_fd_sc_hd__inv_2 _08720_ (.A(net565),
    .Y(_03214_));
 sky130_fd_sc_hd__inv_2 _08721_ (.A(net583),
    .Y(_03225_));
 sky130_fd_sc_hd__inv_2 _08722_ (.A(net602),
    .Y(_03236_));
 sky130_fd_sc_hd__inv_2 _08723_ (.A(net612),
    .Y(_03247_));
 sky130_fd_sc_hd__clkinv_4 _08724_ (.A(net628),
    .Y(_03258_));
 sky130_fd_sc_hd__clkinv_4 _08725_ (.A(net805),
    .Y(_03269_));
 sky130_fd_sc_hd__clkinv_4 _08726_ (.A(net899),
    .Y(_03280_));
 sky130_fd_sc_hd__clkinv_2 _08727_ (.A(net908),
    .Y(_03291_));
 sky130_fd_sc_hd__clkinv_8 _08728_ (.A(net916),
    .Y(_03302_));
 sky130_fd_sc_hd__inv_2 _08729_ (.A(net27),
    .Y(_03313_));
 sky130_fd_sc_hd__inv_2 _08730_ (.A(net69),
    .Y(_03324_));
 sky130_fd_sc_hd__clkinv_4 _08731_ (.A(net313),
    .Y(_03335_));
 sky130_fd_sc_hd__and2_1 _08732_ (.A(net316),
    .B(net315),
    .X(_03346_));
 sky130_fd_sc_hd__nand2_2 _08733_ (.A(net316),
    .B(net315),
    .Y(_03357_));
 sky130_fd_sc_hd__and2b_2 _08734_ (.A_N(\op_code[1] ),
    .B(\op_code[0] ),
    .X(_03367_));
 sky130_fd_sc_hd__mux2_1 _08735_ (.A0(net310),
    .A1(_03367_),
    .S(net280),
    .X(_00002_));
 sky130_fd_sc_hd__nand2_4 _08736_ (.A(\op_code[0] ),
    .B(\op_code[1] ),
    .Y(_03388_));
 sky130_fd_sc_hd__inv_2 _08737_ (.A(_03388_),
    .Y(_03399_));
 sky130_fd_sc_hd__mux2_1 _08738_ (.A0(\sel_op[3] ),
    .A1(_03399_),
    .S(net280),
    .X(_00003_));
 sky130_fd_sc_hd__nand2b_4 _08739_ (.A_N(\op_code[0] ),
    .B(\op_code[1] ),
    .Y(_03420_));
 sky130_fd_sc_hd__nor2_1 _08740_ (.A(net277),
    .B(_03420_),
    .Y(_03431_));
 sky130_fd_sc_hd__a21o_1 _08741_ (.A1(net311),
    .A2(net277),
    .B1(_03431_),
    .X(_00001_));
 sky130_fd_sc_hd__or2_4 _08742_ (.A(\op_code[0] ),
    .B(\op_code[1] ),
    .X(_03452_));
 sky130_fd_sc_hd__nor2_1 _08743_ (.A(net277),
    .B(_03452_),
    .Y(_03463_));
 sky130_fd_sc_hd__a21o_1 _08744_ (.A1(net312),
    .A2(net277),
    .B1(_03463_),
    .X(_00000_));
 sky130_fd_sc_hd__a22o_1 _08745_ (.A1(net421),
    .A2(net756),
    .B1(net777),
    .B2(net404),
    .X(_03484_));
 sky130_fd_sc_hd__and4_1 _08746_ (.A(net404),
    .B(net420),
    .C(net756),
    .D(net777),
    .X(_03495_));
 sky130_fd_sc_hd__inv_2 _08747_ (.A(_03495_),
    .Y(_03506_));
 sky130_fd_sc_hd__and2_2 _08748_ (.A(_03484_),
    .B(_03506_),
    .X(_03517_));
 sky130_fd_sc_hd__nand2_2 _08749_ (.A(net413),
    .B(net767),
    .Y(_03528_));
 sky130_fd_sc_hd__xnor2_4 _08750_ (.A(_03517_),
    .B(_03528_),
    .Y(_03538_));
 sky130_fd_sc_hd__and4_1 _08751_ (.A(net403),
    .B(net421),
    .C(net767),
    .D(net788),
    .X(_03549_));
 sky130_fd_sc_hd__inv_2 _08752_ (.A(_03549_),
    .Y(_03560_));
 sky130_fd_sc_hd__a22o_2 _08753_ (.A1(net419),
    .A2(net767),
    .B1(net788),
    .B2(net403),
    .X(_03571_));
 sky130_fd_sc_hd__and4_2 _08754_ (.A(net411),
    .B(net777),
    .C(_03560_),
    .D(_03571_),
    .X(_03582_));
 sky130_fd_sc_hd__nor2_2 _08755_ (.A(_03549_),
    .B(_03582_),
    .Y(_03593_));
 sky130_fd_sc_hd__nand2b_2 _08756_ (.A_N(_03593_),
    .B(_03538_),
    .Y(_03604_));
 sky130_fd_sc_hd__xor2_4 _08757_ (.A(_03538_),
    .B(_03593_),
    .X(_03615_));
 sky130_fd_sc_hd__a22o_1 _08758_ (.A1(net437),
    .A2(net738),
    .B1(net747),
    .B2(net428),
    .X(_03626_));
 sky130_fd_sc_hd__and2_4 _08759_ (.A(net437),
    .B(net746),
    .X(_03637_));
 sky130_fd_sc_hd__nand2_8 _08760_ (.A(net437),
    .B(net747),
    .Y(_03648_));
 sky130_fd_sc_hd__nand2_8 _08761_ (.A(net427),
    .B(net738),
    .Y(_03659_));
 sky130_fd_sc_hd__o21ai_4 _08762_ (.A1(_03648_),
    .A2(_03659_),
    .B1(_03626_),
    .Y(_03670_));
 sky130_fd_sc_hd__nand2_4 _08763_ (.A(net446),
    .B(net730),
    .Y(_03681_));
 sky130_fd_sc_hd__xor2_4 _08764_ (.A(_03670_),
    .B(_03681_),
    .X(_03691_));
 sky130_fd_sc_hd__nand2b_2 _08765_ (.A_N(_03615_),
    .B(_03691_),
    .Y(_03702_));
 sky130_fd_sc_hd__xnor2_4 _08766_ (.A(_03615_),
    .B(_03691_),
    .Y(_03713_));
 sky130_fd_sc_hd__a22oi_4 _08767_ (.A1(net411),
    .A2(net777),
    .B1(_03560_),
    .B2(_03571_),
    .Y(_03724_));
 sky130_fd_sc_hd__nor2_4 _08768_ (.A(_03582_),
    .B(_03724_),
    .Y(_03735_));
 sky130_fd_sc_hd__and4_2 _08769_ (.A(net403),
    .B(net419),
    .C(net777),
    .D(net801),
    .X(_03746_));
 sky130_fd_sc_hd__inv_2 _08770_ (.A(_03746_),
    .Y(_03757_));
 sky130_fd_sc_hd__a22o_2 _08771_ (.A1(net419),
    .A2(net778),
    .B1(net800),
    .B2(net403),
    .X(_03768_));
 sky130_fd_sc_hd__and4_4 _08772_ (.A(net411),
    .B(net788),
    .C(_03757_),
    .D(_03768_),
    .X(_03779_));
 sky130_fd_sc_hd__nor2_4 _08773_ (.A(_03746_),
    .B(_03779_),
    .Y(_03790_));
 sky130_fd_sc_hd__and2b_2 _08774_ (.A_N(_03790_),
    .B(_03735_),
    .X(_03801_));
 sky130_fd_sc_hd__a21oi_2 _08775_ (.A1(net427),
    .A2(net755),
    .B1(_03637_),
    .Y(_03812_));
 sky130_fd_sc_hd__and3_2 _08776_ (.A(net427),
    .B(net755),
    .C(_03637_),
    .X(_03823_));
 sky130_fd_sc_hd__nor2_4 _08777_ (.A(_03812_),
    .B(_03823_),
    .Y(_03834_));
 sky130_fd_sc_hd__nand2_2 _08778_ (.A(net446),
    .B(net737),
    .Y(_03845_));
 sky130_fd_sc_hd__xor2_4 _08779_ (.A(_03834_),
    .B(_03845_),
    .X(_03856_));
 sky130_fd_sc_hd__xnor2_4 _08780_ (.A(_03735_),
    .B(_03790_),
    .Y(_03866_));
 sky130_fd_sc_hd__and2b_1 _08781_ (.A_N(_03856_),
    .B(_03866_),
    .X(_03877_));
 sky130_fd_sc_hd__o21ai_4 _08782_ (.A1(_03801_),
    .A2(_03877_),
    .B1(_03713_),
    .Y(_03888_));
 sky130_fd_sc_hd__or3_4 _08783_ (.A(_03713_),
    .B(_03801_),
    .C(_03877_),
    .X(_03899_));
 sky130_fd_sc_hd__and4_2 _08784_ (.A(net454),
    .B(net464),
    .C(net720),
    .D(net729),
    .X(_03910_));
 sky130_fd_sc_hd__a22o_1 _08785_ (.A1(net464),
    .A2(net721),
    .B1(net729),
    .B2(net454),
    .X(_03921_));
 sky130_fd_sc_hd__inv_2 _08786_ (.A(_03921_),
    .Y(_03932_));
 sky130_fd_sc_hd__and4b_2 _08787_ (.A_N(_03910_),
    .B(_03921_),
    .C(net474),
    .D(net711),
    .X(_03943_));
 sky130_fd_sc_hd__a31o_2 _08788_ (.A1(net446),
    .A2(net737),
    .A3(_03834_),
    .B1(_03823_),
    .X(_03954_));
 sky130_fd_sc_hd__a22o_1 _08789_ (.A1(net464),
    .A2(net712),
    .B1(net720),
    .B2(net454),
    .X(_03965_));
 sky130_fd_sc_hd__inv_2 _08790_ (.A(_03965_),
    .Y(_03976_));
 sky130_fd_sc_hd__and4_1 _08791_ (.A(net454),
    .B(net464),
    .C(net711),
    .D(net720),
    .X(_03987_));
 sky130_fd_sc_hd__and4b_1 _08792_ (.A_N(_03987_),
    .B(net702),
    .C(net474),
    .D(_03965_),
    .X(_03998_));
 sky130_fd_sc_hd__o2bb2a_1 _08793_ (.A1_N(net474),
    .A2_N(net702),
    .B1(_03976_),
    .B2(_03987_),
    .X(_04008_));
 sky130_fd_sc_hd__nor2_2 _08794_ (.A(_03998_),
    .B(_04008_),
    .Y(_04019_));
 sky130_fd_sc_hd__nand2_1 _08795_ (.A(_03954_),
    .B(_04019_),
    .Y(_04030_));
 sky130_fd_sc_hd__xor2_2 _08796_ (.A(_03954_),
    .B(_04019_),
    .X(_04041_));
 sky130_fd_sc_hd__o21ai_2 _08797_ (.A1(_03910_),
    .A2(_03943_),
    .B1(_04041_),
    .Y(_04052_));
 sky130_fd_sc_hd__or3_1 _08798_ (.A(_03910_),
    .B(_03943_),
    .C(_04041_),
    .X(_04063_));
 sky130_fd_sc_hd__and2_2 _08799_ (.A(_04052_),
    .B(_04063_),
    .X(_04074_));
 sky130_fd_sc_hd__a21o_2 _08800_ (.A1(_03888_),
    .A2(_03899_),
    .B1(_04074_),
    .X(_04085_));
 sky130_fd_sc_hd__nand3_4 _08801_ (.A(_03888_),
    .B(_03899_),
    .C(_04074_),
    .Y(_04096_));
 sky130_fd_sc_hd__xnor2_4 _08802_ (.A(_03856_),
    .B(_03866_),
    .Y(_04107_));
 sky130_fd_sc_hd__a22oi_4 _08803_ (.A1(net411),
    .A2(net788),
    .B1(_03757_),
    .B2(_03768_),
    .Y(_04118_));
 sky130_fd_sc_hd__nor2_4 _08804_ (.A(_03779_),
    .B(_04118_),
    .Y(_04129_));
 sky130_fd_sc_hd__and4_2 _08805_ (.A(net403),
    .B(net419),
    .C(net788),
    .D(net811),
    .X(_04140_));
 sky130_fd_sc_hd__a22oi_2 _08806_ (.A1(net419),
    .A2(net788),
    .B1(net811),
    .B2(net403),
    .Y(_04150_));
 sky130_fd_sc_hd__and4bb_4 _08807_ (.A_N(_04140_),
    .B_N(_04150_),
    .C(net411),
    .D(net801),
    .X(_04161_));
 sky130_fd_sc_hd__nor2_4 _08808_ (.A(_04140_),
    .B(_04161_),
    .Y(_04172_));
 sky130_fd_sc_hd__and2b_2 _08809_ (.A_N(_04172_),
    .B(_04129_),
    .X(_04183_));
 sky130_fd_sc_hd__a22oi_4 _08810_ (.A1(net437),
    .A2(net755),
    .B1(net766),
    .B2(net427),
    .Y(_04194_));
 sky130_fd_sc_hd__and4_1 _08811_ (.A(net427),
    .B(net437),
    .C(net755),
    .D(net766),
    .X(_04205_));
 sky130_fd_sc_hd__nor2_2 _08812_ (.A(_04194_),
    .B(_04205_),
    .Y(_04216_));
 sky130_fd_sc_hd__nand2_4 _08813_ (.A(net446),
    .B(net746),
    .Y(_04227_));
 sky130_fd_sc_hd__xnor2_4 _08814_ (.A(_04216_),
    .B(_04227_),
    .Y(_04238_));
 sky130_fd_sc_hd__xnor2_4 _08815_ (.A(_04129_),
    .B(_04172_),
    .Y(_04249_));
 sky130_fd_sc_hd__and2_2 _08816_ (.A(_04238_),
    .B(_04249_),
    .X(_04260_));
 sky130_fd_sc_hd__o21a_4 _08817_ (.A1(_04183_),
    .A2(_04260_),
    .B1(_04107_),
    .X(_04270_));
 sky130_fd_sc_hd__o21ba_1 _08818_ (.A1(_04194_),
    .A2(_04227_),
    .B1_N(_04205_),
    .X(_04281_));
 sky130_fd_sc_hd__o2bb2a_1 _08819_ (.A1_N(net474),
    .A2_N(net711),
    .B1(_03910_),
    .B2(_03932_),
    .X(_04292_));
 sky130_fd_sc_hd__nor2_1 _08820_ (.A(_03943_),
    .B(_04292_),
    .Y(_04303_));
 sky130_fd_sc_hd__or3_2 _08821_ (.A(_03943_),
    .B(_04281_),
    .C(_04292_),
    .X(_04314_));
 sky130_fd_sc_hd__xnor2_1 _08822_ (.A(_04281_),
    .B(_04303_),
    .Y(_04325_));
 sky130_fd_sc_hd__and4_1 _08823_ (.A(net454),
    .B(net464),
    .C(net729),
    .D(net737),
    .X(_04336_));
 sky130_fd_sc_hd__nand2_4 _08824_ (.A(net474),
    .B(net720),
    .Y(_04347_));
 sky130_fd_sc_hd__a22oi_4 _08825_ (.A1(net464),
    .A2(net729),
    .B1(net737),
    .B2(net454),
    .Y(_04358_));
 sky130_fd_sc_hd__nor2_2 _08826_ (.A(_04336_),
    .B(_04358_),
    .Y(_04369_));
 sky130_fd_sc_hd__o21ba_1 _08827_ (.A1(_04347_),
    .A2(_04358_),
    .B1_N(_04336_),
    .X(_04380_));
 sky130_fd_sc_hd__nand2b_1 _08828_ (.A_N(_04325_),
    .B(_04380_),
    .Y(_04391_));
 sky130_fd_sc_hd__nand2b_2 _08829_ (.A_N(_04380_),
    .B(_04325_),
    .Y(_04402_));
 sky130_fd_sc_hd__nand2_2 _08830_ (.A(_04391_),
    .B(_04402_),
    .Y(_04412_));
 sky130_fd_sc_hd__nor3_4 _08831_ (.A(_04107_),
    .B(_04183_),
    .C(_04260_),
    .Y(_04423_));
 sky130_fd_sc_hd__nor3_4 _08832_ (.A(_04270_),
    .B(_04412_),
    .C(_04423_),
    .Y(_04434_));
 sky130_fd_sc_hd__o211a_4 _08833_ (.A1(_04270_),
    .A2(_04434_),
    .B1(_04085_),
    .C1(_04096_),
    .X(_04445_));
 sky130_fd_sc_hd__a211oi_4 _08834_ (.A1(_04085_),
    .A2(_04096_),
    .B1(_04270_),
    .C1(_04434_),
    .Y(_04456_));
 sky130_fd_sc_hd__a22oi_2 _08835_ (.A1(net491),
    .A2(net694),
    .B1(net702),
    .B2(net481),
    .Y(_04467_));
 sky130_fd_sc_hd__and4_1 _08836_ (.A(net481),
    .B(net491),
    .C(net694),
    .D(net702),
    .X(_04478_));
 sky130_fd_sc_hd__and4bb_1 _08837_ (.A_N(_04467_),
    .B_N(_04478_),
    .C(net501),
    .D(net685),
    .X(_04489_));
 sky130_fd_sc_hd__o2bb2a_1 _08838_ (.A1_N(net501),
    .A2_N(net685),
    .B1(_04467_),
    .B2(_04478_),
    .X(_04500_));
 sky130_fd_sc_hd__nor2_1 _08839_ (.A(_04489_),
    .B(_04500_),
    .Y(_04511_));
 sky130_fd_sc_hd__and4_1 _08840_ (.A(net481),
    .B(net491),
    .C(net702),
    .D(net711),
    .X(_04522_));
 sky130_fd_sc_hd__a22oi_2 _08841_ (.A1(net491),
    .A2(net702),
    .B1(net711),
    .B2(net481),
    .Y(_04532_));
 sky130_fd_sc_hd__and4bb_1 _08842_ (.A_N(_04522_),
    .B_N(_04532_),
    .C(net501),
    .D(net694),
    .X(_04543_));
 sky130_fd_sc_hd__nor2_1 _08843_ (.A(_04522_),
    .B(_04543_),
    .Y(_04554_));
 sky130_fd_sc_hd__and2b_2 _08844_ (.A_N(_04554_),
    .B(_04511_),
    .X(_04565_));
 sky130_fd_sc_hd__xnor2_1 _08845_ (.A(_04511_),
    .B(_04554_),
    .Y(_04576_));
 sky130_fd_sc_hd__a22oi_2 _08846_ (.A1(net517),
    .A2(net667),
    .B1(net676),
    .B2(net508),
    .Y(_04587_));
 sky130_fd_sc_hd__and4_2 _08847_ (.A(net508),
    .B(net517),
    .C(net667),
    .D(net676),
    .X(_04598_));
 sky130_fd_sc_hd__and4bb_2 _08848_ (.A_N(_04587_),
    .B_N(_04598_),
    .C(net525),
    .D(net659),
    .X(_04609_));
 sky130_fd_sc_hd__o2bb2a_1 _08849_ (.A1_N(net525),
    .A2_N(net659),
    .B1(_04587_),
    .B2(_04598_),
    .X(_04620_));
 sky130_fd_sc_hd__nor2_1 _08850_ (.A(_04609_),
    .B(_04620_),
    .Y(_04631_));
 sky130_fd_sc_hd__and2_2 _08851_ (.A(_04576_),
    .B(_04631_),
    .X(_04642_));
 sky130_fd_sc_hd__a22oi_1 _08852_ (.A1(net518),
    .A2(net659),
    .B1(net667),
    .B2(net508),
    .Y(_04652_));
 sky130_fd_sc_hd__and4_1 _08853_ (.A(net508),
    .B(net518),
    .C(net659),
    .D(net667),
    .X(_04663_));
 sky130_fd_sc_hd__nor2_1 _08854_ (.A(_04652_),
    .B(_04663_),
    .Y(_04674_));
 sky130_fd_sc_hd__nand2_1 _08855_ (.A(net526),
    .B(net651),
    .Y(_04685_));
 sky130_fd_sc_hd__xnor2_1 _08856_ (.A(_04674_),
    .B(_04685_),
    .Y(_04696_));
 sky130_fd_sc_hd__a22oi_2 _08857_ (.A1(net492),
    .A2(net685),
    .B1(net694),
    .B2(net482),
    .Y(_04707_));
 sky130_fd_sc_hd__and4_1 _08858_ (.A(net482),
    .B(net492),
    .C(net685),
    .D(net694),
    .X(_04718_));
 sky130_fd_sc_hd__nor2_1 _08859_ (.A(_04707_),
    .B(_04718_),
    .Y(_04729_));
 sky130_fd_sc_hd__nand2_2 _08860_ (.A(net502),
    .B(net677),
    .Y(_04740_));
 sky130_fd_sc_hd__xnor2_2 _08861_ (.A(_04729_),
    .B(_04740_),
    .Y(_04751_));
 sky130_fd_sc_hd__nor2_1 _08862_ (.A(_04478_),
    .B(_04489_),
    .Y(_04761_));
 sky130_fd_sc_hd__and2b_2 _08863_ (.A_N(_04761_),
    .B(_04751_),
    .X(_04772_));
 sky130_fd_sc_hd__xnor2_1 _08864_ (.A(_04751_),
    .B(_04761_),
    .Y(_04783_));
 sky130_fd_sc_hd__and2_2 _08865_ (.A(_04696_),
    .B(_04783_),
    .X(_04794_));
 sky130_fd_sc_hd__nor2_1 _08866_ (.A(_04696_),
    .B(_04783_),
    .Y(_04805_));
 sky130_fd_sc_hd__or2_2 _08867_ (.A(_04794_),
    .B(_04805_),
    .X(_04816_));
 sky130_fd_sc_hd__a21o_4 _08868_ (.A1(_04314_),
    .A2(_04402_),
    .B1(_04816_),
    .X(_04827_));
 sky130_fd_sc_hd__nand3_2 _08869_ (.A(_04314_),
    .B(_04402_),
    .C(_04816_),
    .Y(_04838_));
 sky130_fd_sc_hd__o211ai_4 _08870_ (.A1(_04565_),
    .A2(_04642_),
    .B1(_04827_),
    .C1(_04838_),
    .Y(_04849_));
 sky130_fd_sc_hd__a211o_1 _08871_ (.A1(_04827_),
    .A2(_04838_),
    .B1(_04565_),
    .C1(_04642_),
    .X(_04860_));
 sky130_fd_sc_hd__a2bb2o_2 _08872_ (.A1_N(_04445_),
    .A2_N(_04456_),
    .B1(_04849_),
    .B2(_04860_),
    .X(_04871_));
 sky130_fd_sc_hd__and4bb_2 _08873_ (.A_N(_04445_),
    .B_N(_04456_),
    .C(_04849_),
    .D(_04860_),
    .X(_04881_));
 sky130_fd_sc_hd__or4bb_4 _08874_ (.A(_04445_),
    .B(_04456_),
    .C_N(_04849_),
    .D_N(_04860_),
    .X(_04892_));
 sky130_fd_sc_hd__o21a_2 _08875_ (.A1(_04270_),
    .A2(_04423_),
    .B1(_04412_),
    .X(_04903_));
 sky130_fd_sc_hd__xnor2_4 _08876_ (.A(_04238_),
    .B(_04249_),
    .Y(_04914_));
 sky130_fd_sc_hd__o2bb2a_1 _08877_ (.A1_N(net411),
    .A2_N(net801),
    .B1(_04140_),
    .B2(_04150_),
    .X(_04925_));
 sky130_fd_sc_hd__nor2_2 _08878_ (.A(_04161_),
    .B(_04925_),
    .Y(_04936_));
 sky130_fd_sc_hd__and4_2 _08879_ (.A(net403),
    .B(net419),
    .C(net801),
    .D(net822),
    .X(_04947_));
 sky130_fd_sc_hd__a22oi_2 _08880_ (.A1(net419),
    .A2(net800),
    .B1(net822),
    .B2(net403),
    .Y(_04958_));
 sky130_fd_sc_hd__and4bb_4 _08881_ (.A_N(_04947_),
    .B_N(_04958_),
    .C(net411),
    .D(net811),
    .X(_04969_));
 sky130_fd_sc_hd__nor2_4 _08882_ (.A(_04947_),
    .B(_04969_),
    .Y(_04979_));
 sky130_fd_sc_hd__or3_4 _08883_ (.A(_04161_),
    .B(_04925_),
    .C(_04979_),
    .X(_04990_));
 sky130_fd_sc_hd__nand2_8 _08884_ (.A(net451),
    .B(net763),
    .Y(_05001_));
 sky130_fd_sc_hd__a22oi_4 _08885_ (.A1(net437),
    .A2(net766),
    .B1(net777),
    .B2(net427),
    .Y(_05012_));
 sky130_fd_sc_hd__and4_1 _08886_ (.A(net427),
    .B(net437),
    .C(net766),
    .D(net777),
    .X(_05023_));
 sky130_fd_sc_hd__nor2_2 _08887_ (.A(_05012_),
    .B(_05023_),
    .Y(_05034_));
 sky130_fd_sc_hd__xnor2_4 _08888_ (.A(_05001_),
    .B(_05034_),
    .Y(_05045_));
 sky130_fd_sc_hd__xnor2_4 _08889_ (.A(_04936_),
    .B(_04979_),
    .Y(_05056_));
 sky130_fd_sc_hd__nand2_2 _08890_ (.A(_05045_),
    .B(_05056_),
    .Y(_05067_));
 sky130_fd_sc_hd__a21o_4 _08891_ (.A1(_04990_),
    .A2(_05067_),
    .B1(_04914_),
    .X(_05077_));
 sky130_fd_sc_hd__o21ba_4 _08892_ (.A1(_05001_),
    .A2(_05012_),
    .B1_N(_05023_),
    .X(_05088_));
 sky130_fd_sc_hd__xnor2_4 _08893_ (.A(_04347_),
    .B(_04369_),
    .Y(_05099_));
 sky130_fd_sc_hd__nand2b_1 _08894_ (.A_N(_05088_),
    .B(_05099_),
    .Y(_05110_));
 sky130_fd_sc_hd__xnor2_4 _08895_ (.A(_05088_),
    .B(_05099_),
    .Y(_05121_));
 sky130_fd_sc_hd__nand2_1 _08896_ (.A(net464),
    .B(net746),
    .Y(_05132_));
 sky130_fd_sc_hd__and4_1 _08897_ (.A(net463),
    .B(net473),
    .C(net737),
    .D(net746),
    .X(_05143_));
 sky130_fd_sc_hd__nand2_4 _08898_ (.A(net477),
    .B(net729),
    .Y(_05154_));
 sky130_fd_sc_hd__a22oi_4 _08899_ (.A1(net473),
    .A2(net737),
    .B1(net746),
    .B2(net463),
    .Y(_05164_));
 sky130_fd_sc_hd__nor2_2 _08900_ (.A(_05143_),
    .B(_05164_),
    .Y(_05175_));
 sky130_fd_sc_hd__o21ba_2 _08901_ (.A1(_05154_),
    .A2(_05164_),
    .B1_N(_05143_),
    .X(_05186_));
 sky130_fd_sc_hd__nand2b_1 _08902_ (.A_N(_05186_),
    .B(_05121_),
    .Y(_05197_));
 sky130_fd_sc_hd__xnor2_4 _08903_ (.A(_05121_),
    .B(_05186_),
    .Y(_05208_));
 sky130_fd_sc_hd__nand3_4 _08904_ (.A(_04914_),
    .B(_04990_),
    .C(_05067_),
    .Y(_05219_));
 sky130_fd_sc_hd__nand3_4 _08905_ (.A(_05077_),
    .B(_05208_),
    .C(_05219_),
    .Y(_05230_));
 sky130_fd_sc_hd__a211oi_4 _08906_ (.A1(_05077_),
    .A2(_05230_),
    .B1(_04434_),
    .C1(_04903_),
    .Y(_05241_));
 sky130_fd_sc_hd__nor2_1 _08907_ (.A(_04576_),
    .B(_04631_),
    .Y(_05251_));
 sky130_fd_sc_hd__or2_1 _08908_ (.A(_04642_),
    .B(_05251_),
    .X(_05262_));
 sky130_fd_sc_hd__a21o_2 _08909_ (.A1(_05110_),
    .A2(_05197_),
    .B1(_05262_),
    .X(_05273_));
 sky130_fd_sc_hd__nand3_2 _08910_ (.A(_05110_),
    .B(_05197_),
    .C(_05262_),
    .Y(_05284_));
 sky130_fd_sc_hd__o2bb2a_1 _08911_ (.A1_N(net501),
    .A2_N(net694),
    .B1(_04522_),
    .B2(_04532_),
    .X(_05295_));
 sky130_fd_sc_hd__nor2_1 _08912_ (.A(_04543_),
    .B(_05295_),
    .Y(_05306_));
 sky130_fd_sc_hd__and4_1 _08913_ (.A(net481),
    .B(net491),
    .C(net712),
    .D(net720),
    .X(_05317_));
 sky130_fd_sc_hd__a22oi_2 _08914_ (.A1(net491),
    .A2(net711),
    .B1(net720),
    .B2(net481),
    .Y(_05327_));
 sky130_fd_sc_hd__and4bb_1 _08915_ (.A_N(_05317_),
    .B_N(_05327_),
    .C(net501),
    .D(net702),
    .X(_05338_));
 sky130_fd_sc_hd__nor2_1 _08916_ (.A(_05317_),
    .B(_05338_),
    .Y(_05349_));
 sky130_fd_sc_hd__and2b_2 _08917_ (.A_N(_05349_),
    .B(_05306_),
    .X(_05360_));
 sky130_fd_sc_hd__xnor2_1 _08918_ (.A(_05306_),
    .B(_05349_),
    .Y(_05371_));
 sky130_fd_sc_hd__nand2_1 _08919_ (.A(net525),
    .B(net667),
    .Y(_05382_));
 sky130_fd_sc_hd__a22oi_2 _08920_ (.A1(net517),
    .A2(net676),
    .B1(net685),
    .B2(net508),
    .Y(_05393_));
 sky130_fd_sc_hd__and4_1 _08921_ (.A(net508),
    .B(net517),
    .C(net676),
    .D(net685),
    .X(_05403_));
 sky130_fd_sc_hd__nor2_1 _08922_ (.A(_05393_),
    .B(_05403_),
    .Y(_05414_));
 sky130_fd_sc_hd__xnor2_1 _08923_ (.A(_05382_),
    .B(_05414_),
    .Y(_05425_));
 sky130_fd_sc_hd__and2_2 _08924_ (.A(_05371_),
    .B(_05425_),
    .X(_05436_));
 sky130_fd_sc_hd__a211o_1 _08925_ (.A1(_05273_),
    .A2(_05284_),
    .B1(_05360_),
    .C1(_05436_),
    .X(_05447_));
 sky130_fd_sc_hd__o211ai_4 _08926_ (.A1(_05360_),
    .A2(_05436_),
    .B1(_05273_),
    .C1(_05284_),
    .Y(_05458_));
 sky130_fd_sc_hd__nand2_4 _08927_ (.A(_05447_),
    .B(_05458_),
    .Y(_05468_));
 sky130_fd_sc_hd__o211a_4 _08928_ (.A1(_04434_),
    .A2(_04903_),
    .B1(_05077_),
    .C1(_05230_),
    .X(_05479_));
 sky130_fd_sc_hd__nor3_4 _08929_ (.A(net121),
    .B(_05468_),
    .C(_05479_),
    .Y(_05490_));
 sky130_fd_sc_hd__or3_4 _08930_ (.A(net121),
    .B(_05468_),
    .C(_05479_),
    .X(_05501_));
 sky130_fd_sc_hd__o211ai_4 _08931_ (.A1(_05241_),
    .A2(_05490_),
    .B1(_04871_),
    .C1(_04892_),
    .Y(_05512_));
 sky130_fd_sc_hd__a211o_4 _08932_ (.A1(_04871_),
    .A2(_04892_),
    .B1(_05241_),
    .C1(_05490_),
    .X(_05523_));
 sky130_fd_sc_hd__and4_1 _08933_ (.A(net535),
    .B(net550),
    .C(net651),
    .D(net659),
    .X(_05533_));
 sky130_fd_sc_hd__inv_2 _08934_ (.A(_05533_),
    .Y(_05544_));
 sky130_fd_sc_hd__a22o_1 _08935_ (.A1(net550),
    .A2(net651),
    .B1(net659),
    .B2(net535),
    .X(_05555_));
 sky130_fd_sc_hd__and4_1 _08936_ (.A(net564),
    .B(net642),
    .C(_05544_),
    .D(_05555_),
    .X(_05566_));
 sky130_fd_sc_hd__or2_2 _08937_ (.A(_05533_),
    .B(_05566_),
    .X(_05576_));
 sky130_fd_sc_hd__o21ba_2 _08938_ (.A1(_05382_),
    .A2(_05393_),
    .B1_N(_05403_),
    .X(_05587_));
 sky130_fd_sc_hd__a22oi_2 _08939_ (.A1(net550),
    .A2(net642),
    .B1(net651),
    .B2(net535),
    .Y(_05598_));
 sky130_fd_sc_hd__and4_1 _08940_ (.A(net535),
    .B(net550),
    .C(net642),
    .D(net651),
    .X(_05609_));
 sky130_fd_sc_hd__nor2_2 _08941_ (.A(_05598_),
    .B(_05609_),
    .Y(_05620_));
 sky130_fd_sc_hd__nand2_1 _08942_ (.A(net564),
    .B(net633),
    .Y(_05630_));
 sky130_fd_sc_hd__xnor2_2 _08943_ (.A(_05620_),
    .B(_05630_),
    .Y(_05641_));
 sky130_fd_sc_hd__and2b_1 _08944_ (.A_N(_05587_),
    .B(_05641_),
    .X(_05652_));
 sky130_fd_sc_hd__xnor2_2 _08945_ (.A(_05587_),
    .B(_05641_),
    .Y(_05662_));
 sky130_fd_sc_hd__xnor2_1 _08946_ (.A(_05576_),
    .B(_05662_),
    .Y(_05673_));
 sky130_fd_sc_hd__and4_1 _08947_ (.A(net508),
    .B(net517),
    .C(net685),
    .D(net694),
    .X(_05684_));
 sky130_fd_sc_hd__a22oi_2 _08948_ (.A1(net517),
    .A2(net685),
    .B1(net694),
    .B2(net508),
    .Y(_05695_));
 sky130_fd_sc_hd__and4bb_1 _08949_ (.A_N(_05684_),
    .B_N(_05695_),
    .C(net525),
    .D(net676),
    .X(_05705_));
 sky130_fd_sc_hd__nor2_2 _08950_ (.A(_05684_),
    .B(_05705_),
    .Y(_05716_));
 sky130_fd_sc_hd__a22oi_2 _08951_ (.A1(net564),
    .A2(net642),
    .B1(_05544_),
    .B2(_05555_),
    .Y(_05727_));
 sky130_fd_sc_hd__nor2_1 _08952_ (.A(_05566_),
    .B(_05727_),
    .Y(_05737_));
 sky130_fd_sc_hd__or3_1 _08953_ (.A(_05566_),
    .B(_05716_),
    .C(_05727_),
    .X(_05748_));
 sky130_fd_sc_hd__and4_1 _08954_ (.A(net535),
    .B(net550),
    .C(net659),
    .D(net667),
    .X(_05758_));
 sky130_fd_sc_hd__inv_2 _08955_ (.A(_05758_),
    .Y(_05768_));
 sky130_fd_sc_hd__a22o_1 _08956_ (.A1(net550),
    .A2(net659),
    .B1(net667),
    .B2(net535),
    .X(_05779_));
 sky130_fd_sc_hd__and4_1 _08957_ (.A(net564),
    .B(net651),
    .C(_05768_),
    .D(_05779_),
    .X(_05790_));
 sky130_fd_sc_hd__or2_2 _08958_ (.A(_05758_),
    .B(_05790_),
    .X(_05801_));
 sky130_fd_sc_hd__xnor2_2 _08959_ (.A(_05716_),
    .B(_05737_),
    .Y(_05812_));
 sky130_fd_sc_hd__nand2_1 _08960_ (.A(_05801_),
    .B(_05812_),
    .Y(_05823_));
 sky130_fd_sc_hd__a21oi_1 _08961_ (.A1(_05748_),
    .A2(_05823_),
    .B1(_05673_),
    .Y(_05834_));
 sky130_fd_sc_hd__and3_1 _08962_ (.A(_05673_),
    .B(_05748_),
    .C(_05823_),
    .X(_05845_));
 sky130_fd_sc_hd__a22o_1 _08963_ (.A1(net595),
    .A2(net617),
    .B1(net625),
    .B2(net583),
    .X(_05856_));
 sky130_fd_sc_hd__nand2_4 _08964_ (.A(net595),
    .B(net625),
    .Y(_05867_));
 sky130_fd_sc_hd__nand2_1 _08965_ (.A(net583),
    .B(net617),
    .Y(_05878_));
 sky130_fd_sc_hd__o21a_1 _08966_ (.A1(_05867_),
    .A2(_05878_),
    .B1(_05856_),
    .X(_05888_));
 sky130_fd_sc_hd__and2_4 _08967_ (.A(net606),
    .B(net618),
    .X(_05899_));
 sky130_fd_sc_hd__and2_4 _08968_ (.A(net606),
    .B(net634),
    .X(_05910_));
 sky130_fd_sc_hd__and3_4 _08969_ (.A(net583),
    .B(net617),
    .C(_05910_),
    .X(_05921_));
 sky130_fd_sc_hd__a21oi_4 _08970_ (.A1(net583),
    .A2(net633),
    .B1(_05899_),
    .Y(_05932_));
 sky130_fd_sc_hd__nor3_4 _08971_ (.A(_05867_),
    .B(_05921_),
    .C(_05932_),
    .Y(_05943_));
 sky130_fd_sc_hd__o21ai_4 _08972_ (.A1(_05921_),
    .A2(_05943_),
    .B1(_05888_),
    .Y(_05954_));
 sky130_fd_sc_hd__or3_1 _08973_ (.A(_05888_),
    .B(_05921_),
    .C(_05943_),
    .X(_05965_));
 sky130_fd_sc_hd__and2_1 _08974_ (.A(_05954_),
    .B(_05965_),
    .X(_05976_));
 sky130_fd_sc_hd__a22oi_1 _08975_ (.A1(net326),
    .A2(net892),
    .B1(net901),
    .B2(net317),
    .Y(_05986_));
 sky130_fd_sc_hd__and4_1 _08976_ (.A(net317),
    .B(net326),
    .C(net892),
    .D(net901),
    .X(_05997_));
 sky130_fd_sc_hd__nor2_1 _08977_ (.A(_05986_),
    .B(_05997_),
    .Y(_06008_));
 sky130_fd_sc_hd__and3_1 _08978_ (.A(net335),
    .B(net880),
    .C(_06008_),
    .X(_06019_));
 sky130_fd_sc_hd__a21oi_1 _08979_ (.A1(net335),
    .A2(net880),
    .B1(_06008_),
    .Y(_06030_));
 sky130_fd_sc_hd__or2_1 _08980_ (.A(_06019_),
    .B(_06030_),
    .X(_06040_));
 sky130_fd_sc_hd__inv_2 _08981_ (.A(_06040_),
    .Y(_06051_));
 sky130_fd_sc_hd__nand2_1 _08982_ (.A(_05976_),
    .B(_06051_),
    .Y(_06062_));
 sky130_fd_sc_hd__or2_1 _08983_ (.A(_05976_),
    .B(_06051_),
    .X(_06073_));
 sky130_fd_sc_hd__nand2_1 _08984_ (.A(_06062_),
    .B(_06073_),
    .Y(_06084_));
 sky130_fd_sc_hd__or3_1 _08985_ (.A(_05834_),
    .B(_05845_),
    .C(_06084_),
    .X(_06094_));
 sky130_fd_sc_hd__and2b_2 _08986_ (.A_N(_05834_),
    .B(_06094_),
    .X(_06105_));
 sky130_fd_sc_hd__a22oi_4 _08987_ (.A1(net326),
    .A2(net880),
    .B1(net893),
    .B2(net317),
    .Y(_06116_));
 sky130_fd_sc_hd__and4_1 _08988_ (.A(net317),
    .B(net326),
    .C(net880),
    .D(net892),
    .X(_06127_));
 sky130_fd_sc_hd__nor2_2 _08989_ (.A(_06116_),
    .B(_06127_),
    .Y(_06138_));
 sky130_fd_sc_hd__nand2_4 _08990_ (.A(net335),
    .B(net870),
    .Y(_06149_));
 sky130_fd_sc_hd__xnor2_4 _08991_ (.A(_06138_),
    .B(_06149_),
    .Y(_06160_));
 sky130_fd_sc_hd__inv_2 _08992_ (.A(_06160_),
    .Y(_06170_));
 sky130_fd_sc_hd__and3_1 _08993_ (.A(net583),
    .B(net617),
    .C(_05867_),
    .X(_06181_));
 sky130_fd_sc_hd__xnor2_2 _08994_ (.A(_06160_),
    .B(_06181_),
    .Y(_06192_));
 sky130_fd_sc_hd__a31o_2 _08995_ (.A1(net564),
    .A2(net633),
    .A3(_05620_),
    .B1(_05609_),
    .X(_06203_));
 sky130_fd_sc_hd__nor2_4 _08996_ (.A(_04598_),
    .B(_04609_),
    .Y(_06214_));
 sky130_fd_sc_hd__a22oi_4 _08997_ (.A1(net550),
    .A2(net633),
    .B1(net642),
    .B2(net535),
    .Y(_06225_));
 sky130_fd_sc_hd__and4_2 _08998_ (.A(net535),
    .B(net550),
    .C(net633),
    .D(net642),
    .X(_06235_));
 sky130_fd_sc_hd__nor2_4 _08999_ (.A(_06225_),
    .B(_06235_),
    .Y(_06246_));
 sky130_fd_sc_hd__nand2_2 _09000_ (.A(net564),
    .B(net625),
    .Y(_06257_));
 sky130_fd_sc_hd__xnor2_4 _09001_ (.A(_06246_),
    .B(_06257_),
    .Y(_06268_));
 sky130_fd_sc_hd__and2b_1 _09002_ (.A_N(_06214_),
    .B(_06268_),
    .X(_06279_));
 sky130_fd_sc_hd__xnor2_4 _09003_ (.A(_06214_),
    .B(_06268_),
    .Y(_06290_));
 sky130_fd_sc_hd__xnor2_2 _09004_ (.A(_06203_),
    .B(_06290_),
    .Y(_06301_));
 sky130_fd_sc_hd__a21oi_2 _09005_ (.A1(_05576_),
    .A2(_05662_),
    .B1(_05652_),
    .Y(_06311_));
 sky130_fd_sc_hd__or2_2 _09006_ (.A(_06301_),
    .B(_06311_),
    .X(_06322_));
 sky130_fd_sc_hd__xnor2_1 _09007_ (.A(_06301_),
    .B(_06311_),
    .Y(_06333_));
 sky130_fd_sc_hd__or2_4 _09008_ (.A(_06192_),
    .B(_06333_),
    .X(_06344_));
 sky130_fd_sc_hd__nand2_1 _09009_ (.A(_06192_),
    .B(_06333_),
    .Y(_06355_));
 sky130_fd_sc_hd__nand2_1 _09010_ (.A(_06344_),
    .B(_06355_),
    .Y(_06366_));
 sky130_fd_sc_hd__a21oi_2 _09011_ (.A1(_05273_),
    .A2(_05458_),
    .B1(_06366_),
    .Y(_06376_));
 sky130_fd_sc_hd__and3_1 _09012_ (.A(_05273_),
    .B(_05458_),
    .C(_06366_),
    .X(_06387_));
 sky130_fd_sc_hd__nor2_2 _09013_ (.A(_06376_),
    .B(_06387_),
    .Y(_06398_));
 sky130_fd_sc_hd__xnor2_4 _09014_ (.A(_06105_),
    .B(_06398_),
    .Y(_06409_));
 sky130_fd_sc_hd__and3_2 _09015_ (.A(_05512_),
    .B(_05523_),
    .C(_06409_),
    .X(_06420_));
 sky130_fd_sc_hd__nand3_4 _09016_ (.A(_05512_),
    .B(_05523_),
    .C(_06409_),
    .Y(_06431_));
 sky130_fd_sc_hd__a21oi_4 _09017_ (.A1(_05512_),
    .A2(_05523_),
    .B1(_06409_),
    .Y(_06442_));
 sky130_fd_sc_hd__o21ai_4 _09018_ (.A1(net121),
    .A2(_05479_),
    .B1(_05468_),
    .Y(_06452_));
 sky130_fd_sc_hd__a21o_2 _09019_ (.A1(_05077_),
    .A2(_05219_),
    .B1(_05208_),
    .X(_06463_));
 sky130_fd_sc_hd__xnor2_4 _09020_ (.A(_05045_),
    .B(_05056_),
    .Y(_06474_));
 sky130_fd_sc_hd__o2bb2a_1 _09021_ (.A1_N(net411),
    .A2_N(net811),
    .B1(_04947_),
    .B2(_04958_),
    .X(_06485_));
 sky130_fd_sc_hd__nor2_2 _09022_ (.A(_04969_),
    .B(_06485_),
    .Y(_06496_));
 sky130_fd_sc_hd__and4_2 _09023_ (.A(net403),
    .B(net420),
    .C(net813),
    .D(net831),
    .X(_06507_));
 sky130_fd_sc_hd__a22oi_2 _09024_ (.A1(net420),
    .A2(net813),
    .B1(net832),
    .B2(net405),
    .Y(_06518_));
 sky130_fd_sc_hd__and4bb_4 _09025_ (.A_N(_06507_),
    .B_N(_06518_),
    .C(net411),
    .D(net824),
    .X(_06528_));
 sky130_fd_sc_hd__nor2_4 _09026_ (.A(_06507_),
    .B(_06528_),
    .Y(_06539_));
 sky130_fd_sc_hd__or3_4 _09027_ (.A(_04969_),
    .B(_06485_),
    .C(_06539_),
    .X(_06550_));
 sky130_fd_sc_hd__nand2_8 _09028_ (.A(net448),
    .B(net771),
    .Y(_06561_));
 sky130_fd_sc_hd__a22oi_4 _09029_ (.A1(net436),
    .A2(net777),
    .B1(net788),
    .B2(net427),
    .Y(_06572_));
 sky130_fd_sc_hd__and4_1 _09030_ (.A(net427),
    .B(net436),
    .C(net777),
    .D(net789),
    .X(_06583_));
 sky130_fd_sc_hd__nor2_2 _09031_ (.A(_06572_),
    .B(_06583_),
    .Y(_06594_));
 sky130_fd_sc_hd__xnor2_4 _09032_ (.A(_06561_),
    .B(_06594_),
    .Y(_06605_));
 sky130_fd_sc_hd__xnor2_4 _09033_ (.A(_06496_),
    .B(_06539_),
    .Y(_06615_));
 sky130_fd_sc_hd__nand2_2 _09034_ (.A(_06605_),
    .B(_06615_),
    .Y(_06626_));
 sky130_fd_sc_hd__a21o_2 _09035_ (.A1(_06550_),
    .A2(_06626_),
    .B1(_06474_),
    .X(_06637_));
 sky130_fd_sc_hd__o21ba_4 _09036_ (.A1(_06561_),
    .A2(_06572_),
    .B1_N(_06583_),
    .X(_06648_));
 sky130_fd_sc_hd__xnor2_4 _09037_ (.A(_05154_),
    .B(_05175_),
    .Y(_06659_));
 sky130_fd_sc_hd__nand2b_2 _09038_ (.A_N(_06648_),
    .B(_06659_),
    .Y(_06670_));
 sky130_fd_sc_hd__xnor2_4 _09039_ (.A(_06648_),
    .B(_06659_),
    .Y(_06681_));
 sky130_fd_sc_hd__nand2_8 _09040_ (.A(net458),
    .B(net759),
    .Y(_06692_));
 sky130_fd_sc_hd__nor2_2 _09041_ (.A(_05132_),
    .B(_06692_),
    .Y(_06703_));
 sky130_fd_sc_hd__nand2_2 _09042_ (.A(net474),
    .B(net739),
    .Y(_06713_));
 sky130_fd_sc_hd__nand2_2 _09043_ (.A(_05132_),
    .B(_06692_),
    .Y(_06724_));
 sky130_fd_sc_hd__and2b_2 _09044_ (.A_N(_06703_),
    .B(_06724_),
    .X(_06735_));
 sky130_fd_sc_hd__a31oi_4 _09045_ (.A1(net474),
    .A2(net739),
    .A3(_06724_),
    .B1(_06703_),
    .Y(_06746_));
 sky130_fd_sc_hd__nand2b_2 _09046_ (.A_N(_06746_),
    .B(_06681_),
    .Y(_06757_));
 sky130_fd_sc_hd__xnor2_4 _09047_ (.A(_06681_),
    .B(_06746_),
    .Y(_06768_));
 sky130_fd_sc_hd__nand3_4 _09048_ (.A(_06474_),
    .B(_06550_),
    .C(_06626_),
    .Y(_06779_));
 sky130_fd_sc_hd__nand3_4 _09049_ (.A(_06637_),
    .B(_06768_),
    .C(_06779_),
    .Y(_06790_));
 sky130_fd_sc_hd__nand2_2 _09050_ (.A(_06637_),
    .B(_06790_),
    .Y(_06801_));
 sky130_fd_sc_hd__and3_4 _09051_ (.A(_05230_),
    .B(_06463_),
    .C(_06801_),
    .X(_06811_));
 sky130_fd_sc_hd__nor2_1 _09052_ (.A(_05371_),
    .B(_05425_),
    .Y(_06822_));
 sky130_fd_sc_hd__or2_2 _09053_ (.A(_05436_),
    .B(_06822_),
    .X(_06833_));
 sky130_fd_sc_hd__a21o_4 _09054_ (.A1(_06670_),
    .A2(_06757_),
    .B1(_06833_),
    .X(_06844_));
 sky130_fd_sc_hd__nand3_2 _09055_ (.A(_06670_),
    .B(_06757_),
    .C(_06833_),
    .Y(_06855_));
 sky130_fd_sc_hd__o2bb2a_1 _09056_ (.A1_N(net501),
    .A2_N(net702),
    .B1(_05317_),
    .B2(_05327_),
    .X(_06866_));
 sky130_fd_sc_hd__nor2_1 _09057_ (.A(_05338_),
    .B(_06866_),
    .Y(_06877_));
 sky130_fd_sc_hd__and4_1 _09058_ (.A(net481),
    .B(net491),
    .C(net720),
    .D(net729),
    .X(_06888_));
 sky130_fd_sc_hd__a22oi_2 _09059_ (.A1(net491),
    .A2(net720),
    .B1(net729),
    .B2(net481),
    .Y(_06899_));
 sky130_fd_sc_hd__and4bb_1 _09060_ (.A_N(_06888_),
    .B_N(_06899_),
    .C(net501),
    .D(net711),
    .X(_06909_));
 sky130_fd_sc_hd__nor2_1 _09061_ (.A(_06888_),
    .B(_06909_),
    .Y(_06920_));
 sky130_fd_sc_hd__and2b_2 _09062_ (.A_N(_06920_),
    .B(_06877_),
    .X(_06931_));
 sky130_fd_sc_hd__xnor2_1 _09063_ (.A(_06877_),
    .B(_06920_),
    .Y(_06942_));
 sky130_fd_sc_hd__o2bb2a_1 _09064_ (.A1_N(net525),
    .A2_N(net676),
    .B1(_05684_),
    .B2(_05695_),
    .X(_06953_));
 sky130_fd_sc_hd__nor2_1 _09065_ (.A(_05705_),
    .B(_06953_),
    .Y(_06964_));
 sky130_fd_sc_hd__and2_2 _09066_ (.A(_06942_),
    .B(_06964_),
    .X(_06975_));
 sky130_fd_sc_hd__a211o_1 _09067_ (.A1(_06844_),
    .A2(_06855_),
    .B1(_06931_),
    .C1(_06975_),
    .X(_06986_));
 sky130_fd_sc_hd__o211ai_4 _09068_ (.A1(_06931_),
    .A2(_06975_),
    .B1(_06844_),
    .C1(_06855_),
    .Y(_06997_));
 sky130_fd_sc_hd__nand2_2 _09069_ (.A(_06986_),
    .B(_06997_),
    .Y(_07007_));
 sky130_fd_sc_hd__a21oi_4 _09070_ (.A1(_05230_),
    .A2(_06463_),
    .B1(_06801_),
    .Y(_07018_));
 sky130_fd_sc_hd__nor3_4 _09071_ (.A(_06811_),
    .B(_07007_),
    .C(_07018_),
    .Y(_07029_));
 sky130_fd_sc_hd__o211ai_4 _09072_ (.A1(_06811_),
    .A2(_07029_),
    .B1(_05501_),
    .C1(_06452_),
    .Y(_07040_));
 sky130_fd_sc_hd__o21ai_1 _09073_ (.A1(_05834_),
    .A2(_05845_),
    .B1(_06084_),
    .Y(_07051_));
 sky130_fd_sc_hd__nand2_2 _09074_ (.A(_06094_),
    .B(_07051_),
    .Y(_07062_));
 sky130_fd_sc_hd__a21oi_4 _09075_ (.A1(_06844_),
    .A2(_06997_),
    .B1(_07062_),
    .Y(_07073_));
 sky130_fd_sc_hd__and3_4 _09076_ (.A(_06844_),
    .B(_06997_),
    .C(_07062_),
    .X(_07084_));
 sky130_fd_sc_hd__xnor2_1 _09077_ (.A(_05801_),
    .B(_05812_),
    .Y(_07095_));
 sky130_fd_sc_hd__and4_1 _09078_ (.A(net508),
    .B(net517),
    .C(net695),
    .D(net703),
    .X(_07106_));
 sky130_fd_sc_hd__a22oi_2 _09079_ (.A1(net517),
    .A2(net695),
    .B1(net703),
    .B2(net509),
    .Y(_07117_));
 sky130_fd_sc_hd__and4bb_1 _09080_ (.A_N(_07106_),
    .B_N(_07117_),
    .C(net525),
    .D(net686),
    .X(_07127_));
 sky130_fd_sc_hd__nor2_1 _09081_ (.A(_07106_),
    .B(_07127_),
    .Y(_07138_));
 sky130_fd_sc_hd__a22oi_2 _09082_ (.A1(net564),
    .A2(net652),
    .B1(_05768_),
    .B2(_05779_),
    .Y(_07149_));
 sky130_fd_sc_hd__nor2_1 _09083_ (.A(_05790_),
    .B(_07149_),
    .Y(_07160_));
 sky130_fd_sc_hd__or3_1 _09084_ (.A(_05790_),
    .B(_07138_),
    .C(_07149_),
    .X(_07171_));
 sky130_fd_sc_hd__and4_2 _09085_ (.A(net535),
    .B(net550),
    .C(net667),
    .D(net676),
    .X(_07182_));
 sky130_fd_sc_hd__a22oi_2 _09086_ (.A1(net550),
    .A2(net667),
    .B1(net676),
    .B2(net535),
    .Y(_07193_));
 sky130_fd_sc_hd__and4bb_2 _09087_ (.A_N(_07182_),
    .B_N(_07193_),
    .C(net564),
    .D(net660),
    .X(_07204_));
 sky130_fd_sc_hd__xnor2_1 _09088_ (.A(_07138_),
    .B(_07160_),
    .Y(_07215_));
 sky130_fd_sc_hd__o21ai_2 _09089_ (.A1(_07182_),
    .A2(_07204_),
    .B1(_07215_),
    .Y(_07226_));
 sky130_fd_sc_hd__a21o_1 _09090_ (.A1(_07171_),
    .A2(_07226_),
    .B1(_07095_),
    .X(_07237_));
 sky130_fd_sc_hd__and3_1 _09091_ (.A(_07095_),
    .B(_07171_),
    .C(_07226_),
    .X(_07247_));
 sky130_fd_sc_hd__inv_2 _09092_ (.A(_07247_),
    .Y(_07258_));
 sky130_fd_sc_hd__nand2_2 _09093_ (.A(_07237_),
    .B(_07258_),
    .Y(_07269_));
 sky130_fd_sc_hd__o21a_1 _09094_ (.A1(_05921_),
    .A2(_05932_),
    .B1(_05867_),
    .X(_07280_));
 sky130_fd_sc_hd__nor2_1 _09095_ (.A(_05943_),
    .B(_07280_),
    .Y(_07291_));
 sky130_fd_sc_hd__and2_2 _09096_ (.A(net606),
    .B(net643),
    .X(_07302_));
 sky130_fd_sc_hd__and2_1 _09097_ (.A(net606),
    .B(net626),
    .X(_07313_));
 sky130_fd_sc_hd__and3_1 _09098_ (.A(net583),
    .B(net626),
    .C(_07302_),
    .X(_07324_));
 sky130_fd_sc_hd__a21oi_2 _09099_ (.A1(net583),
    .A2(net643),
    .B1(_07313_),
    .Y(_07335_));
 sky130_fd_sc_hd__and4bb_2 _09100_ (.A_N(_07324_),
    .B_N(_07335_),
    .C(net595),
    .D(net634),
    .X(_07346_));
 sky130_fd_sc_hd__nor2_2 _09101_ (.A(_07324_),
    .B(_07346_),
    .Y(_07356_));
 sky130_fd_sc_hd__and2b_2 _09102_ (.A_N(_07356_),
    .B(_07291_),
    .X(_07367_));
 sky130_fd_sc_hd__xnor2_1 _09103_ (.A(_07291_),
    .B(_07356_),
    .Y(_07378_));
 sky130_fd_sc_hd__a22oi_4 _09104_ (.A1(net326),
    .A2(net901),
    .B1(net910),
    .B2(net317),
    .Y(_07389_));
 sky130_fd_sc_hd__and4_1 _09105_ (.A(net317),
    .B(net326),
    .C(net901),
    .D(net910),
    .X(_07400_));
 sky130_fd_sc_hd__nor2_1 _09106_ (.A(_07389_),
    .B(_07400_),
    .Y(_07411_));
 sky130_fd_sc_hd__nand2_1 _09107_ (.A(net335),
    .B(net892),
    .Y(_07422_));
 sky130_fd_sc_hd__xnor2_1 _09108_ (.A(_07411_),
    .B(_07422_),
    .Y(_07433_));
 sky130_fd_sc_hd__and2_2 _09109_ (.A(_07378_),
    .B(_07433_),
    .X(_07444_));
 sky130_fd_sc_hd__nor2_1 _09110_ (.A(_07378_),
    .B(_07433_),
    .Y(_07454_));
 sky130_fd_sc_hd__or2_4 _09111_ (.A(_07444_),
    .B(_07454_),
    .X(_07465_));
 sky130_fd_sc_hd__o21a_4 _09112_ (.A1(_07247_),
    .A2(_07465_),
    .B1(_07237_),
    .X(_07476_));
 sky130_fd_sc_hd__o21ai_4 _09113_ (.A1(_07073_),
    .A2(_07084_),
    .B1(_07476_),
    .Y(_07487_));
 sky130_fd_sc_hd__nor3_4 _09114_ (.A(_07073_),
    .B(_07084_),
    .C(_07476_),
    .Y(_07498_));
 sky130_fd_sc_hd__or3_4 _09115_ (.A(_07073_),
    .B(_07084_),
    .C(_07476_),
    .X(_07509_));
 sky130_fd_sc_hd__nand2_2 _09116_ (.A(_07487_),
    .B(_07509_),
    .Y(_07520_));
 sky130_fd_sc_hd__a211o_4 _09117_ (.A1(_05501_),
    .A2(_06452_),
    .B1(_06811_),
    .C1(_07029_),
    .X(_07531_));
 sky130_fd_sc_hd__nand2_2 _09118_ (.A(_07040_),
    .B(_07531_),
    .Y(_07542_));
 sky130_fd_sc_hd__nand4_4 _09119_ (.A(_07040_),
    .B(_07487_),
    .C(_07509_),
    .D(_07531_),
    .Y(_07552_));
 sky130_fd_sc_hd__a211oi_4 _09120_ (.A1(_07040_),
    .A2(_07552_),
    .B1(_06420_),
    .C1(_06442_),
    .Y(_07563_));
 sky130_fd_sc_hd__o211a_1 _09121_ (.A1(_06420_),
    .A2(_06442_),
    .B1(_07040_),
    .C1(_07552_),
    .X(_07574_));
 sky130_fd_sc_hd__nor2_4 _09122_ (.A(_07563_),
    .B(_07574_),
    .Y(_07585_));
 sky130_fd_sc_hd__nand2_4 _09123_ (.A(net335),
    .B(net910),
    .Y(_07596_));
 sky130_fd_sc_hd__and4_4 _09124_ (.A(net326),
    .B(net335),
    .C(net901),
    .D(net910),
    .X(_07607_));
 sky130_fd_sc_hd__a22o_1 _09125_ (.A1(net349),
    .A2(net870),
    .B1(net880),
    .B2(net340),
    .X(_07618_));
 sky130_fd_sc_hd__inv_2 _09126_ (.A(_07618_),
    .Y(_07629_));
 sky130_fd_sc_hd__and4_2 _09127_ (.A(net340),
    .B(net349),
    .C(net870),
    .D(net880),
    .X(_07640_));
 sky130_fd_sc_hd__and4b_4 _09128_ (.A_N(_07640_),
    .B(net860),
    .C(net357),
    .D(_07618_),
    .X(_07650_));
 sky130_fd_sc_hd__o2bb2a_1 _09129_ (.A1_N(net357),
    .A2_N(net860),
    .B1(_07629_),
    .B2(_07640_),
    .X(_07661_));
 sky130_fd_sc_hd__nor2_4 _09130_ (.A(_07650_),
    .B(_07661_),
    .Y(_07672_));
 sky130_fd_sc_hd__and2_1 _09131_ (.A(_07607_),
    .B(_07672_),
    .X(_07683_));
 sky130_fd_sc_hd__and4_1 _09132_ (.A(net340),
    .B(net350),
    .C(net880),
    .D(net892),
    .X(_07694_));
 sky130_fd_sc_hd__nand2_1 _09133_ (.A(net357),
    .B(net870),
    .Y(_07705_));
 sky130_fd_sc_hd__a22oi_1 _09134_ (.A1(net350),
    .A2(net880),
    .B1(net892),
    .B2(net340),
    .Y(_07716_));
 sky130_fd_sc_hd__nor2_1 _09135_ (.A(_07694_),
    .B(_07716_),
    .Y(_07727_));
 sky130_fd_sc_hd__a31o_4 _09136_ (.A1(net357),
    .A2(net870),
    .A3(_07727_),
    .B1(_07694_),
    .X(_07738_));
 sky130_fd_sc_hd__xnor2_4 _09137_ (.A(_07607_),
    .B(_07672_),
    .Y(_07748_));
 sky130_fd_sc_hd__and2b_1 _09138_ (.A_N(_07748_),
    .B(_07738_),
    .X(_07759_));
 sky130_fd_sc_hd__nor2_4 _09139_ (.A(_07640_),
    .B(_07650_),
    .Y(_07770_));
 sky130_fd_sc_hd__o21ba_4 _09140_ (.A1(_07389_),
    .A2(_07422_),
    .B1_N(_07400_),
    .X(_07781_));
 sky130_fd_sc_hd__a22oi_1 _09141_ (.A1(net349),
    .A2(net860),
    .B1(net870),
    .B2(net340),
    .Y(_07792_));
 sky130_fd_sc_hd__and4_1 _09142_ (.A(net340),
    .B(net349),
    .C(net860),
    .D(net870),
    .X(_07803_));
 sky130_fd_sc_hd__nor2_1 _09143_ (.A(_07792_),
    .B(_07803_),
    .Y(_07814_));
 sky130_fd_sc_hd__a21oi_1 _09144_ (.A1(net357),
    .A2(net850),
    .B1(_07814_),
    .Y(_07825_));
 sky130_fd_sc_hd__and3_1 _09145_ (.A(net357),
    .B(net850),
    .C(_07814_),
    .X(_07835_));
 sky130_fd_sc_hd__nor2_2 _09146_ (.A(_07825_),
    .B(_07835_),
    .Y(_07846_));
 sky130_fd_sc_hd__or3_2 _09147_ (.A(_07781_),
    .B(_07825_),
    .C(_07835_),
    .X(_07857_));
 sky130_fd_sc_hd__xnor2_4 _09148_ (.A(_07781_),
    .B(_07846_),
    .Y(_07868_));
 sky130_fd_sc_hd__nand2b_2 _09149_ (.A_N(_07770_),
    .B(_07868_),
    .Y(_07879_));
 sky130_fd_sc_hd__xnor2_4 _09150_ (.A(_07770_),
    .B(_07868_),
    .Y(_07890_));
 sky130_fd_sc_hd__o21ai_4 _09151_ (.A1(_07367_),
    .A2(_07444_),
    .B1(_07890_),
    .Y(_07901_));
 sky130_fd_sc_hd__inv_2 _09152_ (.A(_07901_),
    .Y(_07912_));
 sky130_fd_sc_hd__or3_1 _09153_ (.A(_07367_),
    .B(_07444_),
    .C(_07890_),
    .X(_07922_));
 sky130_fd_sc_hd__o211a_2 _09154_ (.A1(_07683_),
    .A2(_07759_),
    .B1(_07901_),
    .C1(_07922_),
    .X(_07933_));
 sky130_fd_sc_hd__inv_2 _09155_ (.A(_07933_),
    .Y(_07944_));
 sky130_fd_sc_hd__a211o_2 _09156_ (.A1(_07901_),
    .A2(_07922_),
    .B1(_07683_),
    .C1(_07759_),
    .X(_07955_));
 sky130_fd_sc_hd__o2bb2a_1 _09157_ (.A1_N(net595),
    .A2_N(net633),
    .B1(_07324_),
    .B2(_07335_),
    .X(_07966_));
 sky130_fd_sc_hd__nor2_2 _09158_ (.A(_07346_),
    .B(_07966_),
    .Y(_07977_));
 sky130_fd_sc_hd__and2_2 _09159_ (.A(net607),
    .B(net653),
    .X(_07987_));
 sky130_fd_sc_hd__and3_2 _09160_ (.A(net581),
    .B(net634),
    .C(_07987_),
    .X(_07998_));
 sky130_fd_sc_hd__inv_2 _09161_ (.A(_07998_),
    .Y(_08009_));
 sky130_fd_sc_hd__a21o_1 _09162_ (.A1(net583),
    .A2(net651),
    .B1(_05910_),
    .X(_08020_));
 sky130_fd_sc_hd__and4b_4 _09163_ (.A_N(_07998_),
    .B(_08020_),
    .C(net595),
    .D(net642),
    .X(_08031_));
 sky130_fd_sc_hd__nor2_4 _09164_ (.A(_07998_),
    .B(_08031_),
    .Y(_08042_));
 sky130_fd_sc_hd__or3_4 _09165_ (.A(_07346_),
    .B(_07966_),
    .C(_08042_),
    .X(_08053_));
 sky130_fd_sc_hd__a22oi_1 _09166_ (.A1(net335),
    .A2(net901),
    .B1(net910),
    .B2(net326),
    .Y(_08063_));
 sky130_fd_sc_hd__or2_4 _09167_ (.A(_07607_),
    .B(_08063_),
    .X(_08074_));
 sky130_fd_sc_hd__xnor2_4 _09168_ (.A(_07977_),
    .B(_08042_),
    .Y(_08085_));
 sky130_fd_sc_hd__nand2b_2 _09169_ (.A_N(_08074_),
    .B(_08085_),
    .Y(_08096_));
 sky130_fd_sc_hd__xor2_4 _09170_ (.A(_07738_),
    .B(_07748_),
    .X(_08107_));
 sky130_fd_sc_hd__a21oi_4 _09171_ (.A1(_08053_),
    .A2(_08096_),
    .B1(_08107_),
    .Y(_08118_));
 sky130_fd_sc_hd__and2_1 _09172_ (.A(net356),
    .B(net901),
    .X(_08128_));
 sky130_fd_sc_hd__and3_1 _09173_ (.A(net341),
    .B(net892),
    .C(_08128_),
    .X(_08139_));
 sky130_fd_sc_hd__a22oi_2 _09174_ (.A1(net356),
    .A2(net892),
    .B1(net901),
    .B2(net341),
    .Y(_08150_));
 sky130_fd_sc_hd__and4bb_1 _09175_ (.A_N(_08139_),
    .B_N(_08150_),
    .C(net358),
    .D(net881),
    .X(_08161_));
 sky130_fd_sc_hd__xnor2_1 _09176_ (.A(_07705_),
    .B(_07727_),
    .Y(_08172_));
 sky130_fd_sc_hd__o21a_1 _09177_ (.A1(_08139_),
    .A2(_08161_),
    .B1(_08172_),
    .X(_08182_));
 sky130_fd_sc_hd__and3_1 _09178_ (.A(_08053_),
    .B(_08096_),
    .C(_08107_),
    .X(_08193_));
 sky130_fd_sc_hd__nor2_1 _09179_ (.A(_08118_),
    .B(_08193_),
    .Y(_08204_));
 sky130_fd_sc_hd__and2_2 _09180_ (.A(_08182_),
    .B(_08204_),
    .X(_08215_));
 sky130_fd_sc_hd__o211ai_4 _09181_ (.A1(_08118_),
    .A2(_08215_),
    .B1(_07944_),
    .C1(_07955_),
    .Y(_08226_));
 sky130_fd_sc_hd__inv_2 _09182_ (.A(_08226_),
    .Y(_08236_));
 sky130_fd_sc_hd__a211o_1 _09183_ (.A1(_07944_),
    .A2(_07955_),
    .B1(_08118_),
    .C1(_08215_),
    .X(_08247_));
 sky130_fd_sc_hd__nand2_1 _09184_ (.A(net396),
    .B(net801),
    .Y(_08258_));
 sky130_fd_sc_hd__a22oi_4 _09185_ (.A1(net372),
    .A2(net830),
    .B1(net840),
    .B2(net363),
    .Y(_08269_));
 sky130_fd_sc_hd__and4_2 _09186_ (.A(net363),
    .B(net372),
    .C(net830),
    .D(net840),
    .X(_08280_));
 sky130_fd_sc_hd__nand2_1 _09187_ (.A(net383),
    .B(net821),
    .Y(_08290_));
 sky130_fd_sc_hd__o21a_1 _09188_ (.A1(_08269_),
    .A2(_08280_),
    .B1(_08290_),
    .X(_08301_));
 sky130_fd_sc_hd__nor3_2 _09189_ (.A(_08269_),
    .B(_08280_),
    .C(_08290_),
    .Y(_08312_));
 sky130_fd_sc_hd__nor2_2 _09190_ (.A(_08301_),
    .B(_08312_),
    .Y(_08322_));
 sky130_fd_sc_hd__and4_2 _09191_ (.A(net363),
    .B(net372),
    .C(net840),
    .D(net850),
    .X(_08333_));
 sky130_fd_sc_hd__a22o_1 _09192_ (.A1(net372),
    .A2(net840),
    .B1(net850),
    .B2(net363),
    .X(_08344_));
 sky130_fd_sc_hd__inv_2 _09193_ (.A(_08344_),
    .Y(_08354_));
 sky130_fd_sc_hd__and4b_2 _09194_ (.A_N(_08333_),
    .B(_08344_),
    .C(net383),
    .D(net830),
    .X(_08365_));
 sky130_fd_sc_hd__o21ai_4 _09195_ (.A1(_08333_),
    .A2(_08365_),
    .B1(_08322_),
    .Y(_08376_));
 sky130_fd_sc_hd__or3_1 _09196_ (.A(_08322_),
    .B(_08333_),
    .C(_08365_),
    .X(_08386_));
 sky130_fd_sc_hd__and2_2 _09197_ (.A(_08376_),
    .B(_08386_),
    .X(_08397_));
 sky130_fd_sc_hd__nand3_4 _09198_ (.A(net388),
    .B(net810),
    .C(_08397_),
    .Y(_08408_));
 sky130_fd_sc_hd__a21o_1 _09199_ (.A1(net388),
    .A2(net810),
    .B1(_08397_),
    .X(_08415_));
 sky130_fd_sc_hd__and2_1 _09200_ (.A(_08408_),
    .B(_08415_),
    .X(_08423_));
 sky130_fd_sc_hd__o2bb2a_1 _09201_ (.A1_N(net383),
    .A2_N(net830),
    .B1(_08333_),
    .B2(_08354_),
    .X(_08431_));
 sky130_fd_sc_hd__nor2_1 _09202_ (.A(_08365_),
    .B(_08431_),
    .Y(_08438_));
 sky130_fd_sc_hd__and4_1 _09203_ (.A(net363),
    .B(net372),
    .C(net851),
    .D(net860),
    .X(_08446_));
 sky130_fd_sc_hd__a22oi_2 _09204_ (.A1(net372),
    .A2(net851),
    .B1(net861),
    .B2(net363),
    .Y(_08454_));
 sky130_fd_sc_hd__and4bb_1 _09205_ (.A_N(_08446_),
    .B_N(_08454_),
    .C(net383),
    .D(net842),
    .X(_08461_));
 sky130_fd_sc_hd__nor2_1 _09206_ (.A(_08446_),
    .B(_08461_),
    .Y(_08469_));
 sky130_fd_sc_hd__and2b_1 _09207_ (.A_N(_08469_),
    .B(_08438_),
    .X(_08477_));
 sky130_fd_sc_hd__xnor2_1 _09208_ (.A(_08438_),
    .B(_08469_),
    .Y(_08485_));
 sky130_fd_sc_hd__and3_2 _09209_ (.A(net388),
    .B(net821),
    .C(_08485_),
    .X(_08491_));
 sky130_fd_sc_hd__o21a_1 _09210_ (.A1(_08477_),
    .A2(_08491_),
    .B1(_08423_),
    .X(_08497_));
 sky130_fd_sc_hd__nor3_1 _09211_ (.A(_08423_),
    .B(_08477_),
    .C(_08491_),
    .Y(_08503_));
 sky130_fd_sc_hd__nor2_2 _09212_ (.A(_08497_),
    .B(_08503_),
    .Y(_08509_));
 sky130_fd_sc_hd__xnor2_1 _09213_ (.A(_08258_),
    .B(_08509_),
    .Y(_08515_));
 sky130_fd_sc_hd__and3_2 _09214_ (.A(_08226_),
    .B(_08247_),
    .C(_08515_),
    .X(_08521_));
 sky130_fd_sc_hd__a22oi_4 _09215_ (.A1(net372),
    .A2(net821),
    .B1(net830),
    .B2(net363),
    .Y(_08528_));
 sky130_fd_sc_hd__and4_2 _09216_ (.A(net363),
    .B(net372),
    .C(net821),
    .D(net830),
    .X(_08534_));
 sky130_fd_sc_hd__nand2_1 _09217_ (.A(net383),
    .B(net810),
    .Y(_08540_));
 sky130_fd_sc_hd__o21a_1 _09218_ (.A1(_08528_),
    .A2(_08534_),
    .B1(_08540_),
    .X(_08546_));
 sky130_fd_sc_hd__nor3_2 _09219_ (.A(_08528_),
    .B(_08534_),
    .C(_08540_),
    .Y(_08552_));
 sky130_fd_sc_hd__nor2_2 _09220_ (.A(_08546_),
    .B(_08552_),
    .Y(_08558_));
 sky130_fd_sc_hd__nor3_2 _09221_ (.A(_08280_),
    .B(_08312_),
    .C(_08558_),
    .Y(_08564_));
 sky130_fd_sc_hd__o21a_2 _09222_ (.A1(_08280_),
    .A2(_08312_),
    .B1(_08558_),
    .X(_08565_));
 sky130_fd_sc_hd__nor2_4 _09223_ (.A(_08564_),
    .B(_08565_),
    .Y(_08566_));
 sky130_fd_sc_hd__nand2_2 _09224_ (.A(net388),
    .B(net800),
    .Y(_08567_));
 sky130_fd_sc_hd__xor2_4 _09225_ (.A(_08566_),
    .B(_08567_),
    .X(_08568_));
 sky130_fd_sc_hd__a21oi_4 _09226_ (.A1(_08376_),
    .A2(_08408_),
    .B1(_08568_),
    .Y(_08569_));
 sky130_fd_sc_hd__and3_1 _09227_ (.A(_08376_),
    .B(_08408_),
    .C(_08568_),
    .X(_08570_));
 sky130_fd_sc_hd__nor2_4 _09228_ (.A(_08569_),
    .B(_08570_),
    .Y(_08571_));
 sky130_fd_sc_hd__nand2_2 _09229_ (.A(net396),
    .B(net790),
    .Y(_08572_));
 sky130_fd_sc_hd__xnor2_4 _09230_ (.A(_08571_),
    .B(_08572_),
    .Y(_08573_));
 sky130_fd_sc_hd__or2_2 _09231_ (.A(_07803_),
    .B(_07835_),
    .X(_08574_));
 sky130_fd_sc_hd__a22oi_2 _09232_ (.A1(net349),
    .A2(net850),
    .B1(net860),
    .B2(net340),
    .Y(_08575_));
 sky130_fd_sc_hd__and4_1 _09233_ (.A(net340),
    .B(net349),
    .C(net850),
    .D(net860),
    .X(_08576_));
 sky130_fd_sc_hd__nor2_1 _09234_ (.A(_08575_),
    .B(_08576_),
    .Y(_08577_));
 sky130_fd_sc_hd__nand2_1 _09235_ (.A(net357),
    .B(net840),
    .Y(_08578_));
 sky130_fd_sc_hd__xnor2_1 _09236_ (.A(_08577_),
    .B(_08578_),
    .Y(_08579_));
 sky130_fd_sc_hd__o21a_1 _09237_ (.A1(_05997_),
    .A2(_06019_),
    .B1(_08579_),
    .X(_08580_));
 sky130_fd_sc_hd__nor3_1 _09238_ (.A(_05997_),
    .B(_06019_),
    .C(_08579_),
    .Y(_08581_));
 sky130_fd_sc_hd__nor2_1 _09239_ (.A(_08580_),
    .B(_08581_),
    .Y(_08582_));
 sky130_fd_sc_hd__xnor2_1 _09240_ (.A(_08574_),
    .B(_08582_),
    .Y(_08583_));
 sky130_fd_sc_hd__a21o_2 _09241_ (.A1(_05954_),
    .A2(_06062_),
    .B1(_08583_),
    .X(_08584_));
 sky130_fd_sc_hd__nand3_1 _09242_ (.A(_05954_),
    .B(_06062_),
    .C(_08583_),
    .Y(_08585_));
 sky130_fd_sc_hd__nand2_2 _09243_ (.A(_08584_),
    .B(_08585_),
    .Y(_08586_));
 sky130_fd_sc_hd__a21o_4 _09244_ (.A1(_07857_),
    .A2(_07879_),
    .B1(_08586_),
    .X(_08587_));
 sky130_fd_sc_hd__nand3_2 _09245_ (.A(_07857_),
    .B(_07879_),
    .C(_08586_),
    .Y(_08588_));
 sky130_fd_sc_hd__o211ai_4 _09246_ (.A1(_07912_),
    .A2(_07933_),
    .B1(_08587_),
    .C1(_08588_),
    .Y(_08589_));
 sky130_fd_sc_hd__a211o_2 _09247_ (.A1(_08587_),
    .A2(_08588_),
    .B1(_07912_),
    .C1(_07933_),
    .X(_08590_));
 sky130_fd_sc_hd__nand3_4 _09248_ (.A(_08573_),
    .B(_08589_),
    .C(_08590_),
    .Y(_08591_));
 sky130_fd_sc_hd__a21o_2 _09249_ (.A1(_08589_),
    .A2(_08590_),
    .B1(_08573_),
    .X(_08592_));
 sky130_fd_sc_hd__o211ai_4 _09250_ (.A1(_07073_),
    .A2(_07498_),
    .B1(_08591_),
    .C1(_08592_),
    .Y(_08593_));
 sky130_fd_sc_hd__a211o_2 _09251_ (.A1(_08591_),
    .A2(_08592_),
    .B1(_07073_),
    .C1(_07498_),
    .X(_08594_));
 sky130_fd_sc_hd__o211ai_4 _09252_ (.A1(_08236_),
    .A2(_08521_),
    .B1(_08593_),
    .C1(_08594_),
    .Y(_08595_));
 sky130_fd_sc_hd__a211o_1 _09253_ (.A1(_08593_),
    .A2(_08594_),
    .B1(_08236_),
    .C1(_08521_),
    .X(_08596_));
 sky130_fd_sc_hd__nand2_2 _09254_ (.A(_08595_),
    .B(_08596_),
    .Y(_08597_));
 sky130_fd_sc_hd__and3_2 _09255_ (.A(_07585_),
    .B(_08595_),
    .C(_08596_),
    .X(_08598_));
 sky130_fd_sc_hd__xnor2_4 _09256_ (.A(_07585_),
    .B(_08597_),
    .Y(_08599_));
 sky130_fd_sc_hd__xnor2_4 _09257_ (.A(_07520_),
    .B(_07542_),
    .Y(_08600_));
 sky130_fd_sc_hd__o21a_1 _09258_ (.A1(_06811_),
    .A2(_07018_),
    .B1(_07007_),
    .X(_08601_));
 sky130_fd_sc_hd__or2_4 _09259_ (.A(_07029_),
    .B(_08601_),
    .X(_08602_));
 sky130_fd_sc_hd__a21o_1 _09260_ (.A1(_06637_),
    .A2(_06779_),
    .B1(_06768_),
    .X(_08603_));
 sky130_fd_sc_hd__nand2_1 _09261_ (.A(_06790_),
    .B(_08603_),
    .Y(_08604_));
 sky130_fd_sc_hd__xnor2_4 _09262_ (.A(_06605_),
    .B(_06615_),
    .Y(_08605_));
 sky130_fd_sc_hd__o2bb2a_1 _09263_ (.A1_N(net411),
    .A2_N(net824),
    .B1(_06507_),
    .B2(_06518_),
    .X(_08606_));
 sky130_fd_sc_hd__nor2_2 _09264_ (.A(_06528_),
    .B(_08606_),
    .Y(_08607_));
 sky130_fd_sc_hd__and4_2 _09265_ (.A(net404),
    .B(net420),
    .C(net824),
    .D(net841),
    .X(_08608_));
 sky130_fd_sc_hd__a22oi_2 _09266_ (.A1(net420),
    .A2(net823),
    .B1(net841),
    .B2(net403),
    .Y(_08609_));
 sky130_fd_sc_hd__and4bb_4 _09267_ (.A_N(_08608_),
    .B_N(_08609_),
    .C(net412),
    .D(net832),
    .X(_08610_));
 sky130_fd_sc_hd__nor2_4 _09268_ (.A(_08608_),
    .B(_08610_),
    .Y(_08611_));
 sky130_fd_sc_hd__or3_4 _09269_ (.A(_06528_),
    .B(_08606_),
    .C(_08611_),
    .X(_08612_));
 sky130_fd_sc_hd__nand2_8 _09270_ (.A(net450),
    .B(net787),
    .Y(_08613_));
 sky130_fd_sc_hd__a22oi_4 _09271_ (.A1(net436),
    .A2(net788),
    .B1(net803),
    .B2(net428),
    .Y(_08614_));
 sky130_fd_sc_hd__and4_1 _09272_ (.A(net427),
    .B(net436),
    .C(net788),
    .D(net803),
    .X(_08615_));
 sky130_fd_sc_hd__nor2_2 _09273_ (.A(_08614_),
    .B(_08615_),
    .Y(_08616_));
 sky130_fd_sc_hd__xnor2_4 _09274_ (.A(_08613_),
    .B(_08616_),
    .Y(_08617_));
 sky130_fd_sc_hd__xnor2_4 _09275_ (.A(_08607_),
    .B(_08611_),
    .Y(_08618_));
 sky130_fd_sc_hd__nand2_2 _09276_ (.A(_08617_),
    .B(_08618_),
    .Y(_08619_));
 sky130_fd_sc_hd__a21o_4 _09277_ (.A1(_08612_),
    .A2(_08619_),
    .B1(_08605_),
    .X(_08620_));
 sky130_fd_sc_hd__o21ba_4 _09278_ (.A1(_08613_),
    .A2(_08614_),
    .B1_N(_08615_),
    .X(_08621_));
 sky130_fd_sc_hd__xnor2_4 _09279_ (.A(_06713_),
    .B(_06735_),
    .Y(_08622_));
 sky130_fd_sc_hd__nand2b_2 _09280_ (.A_N(_08621_),
    .B(_08622_),
    .Y(_08623_));
 sky130_fd_sc_hd__xnor2_4 _09281_ (.A(_08621_),
    .B(_08622_),
    .Y(_08624_));
 sky130_fd_sc_hd__nand2_8 _09282_ (.A(net465),
    .B(net766),
    .Y(_08625_));
 sky130_fd_sc_hd__nand2_8 _09283_ (.A(net458),
    .B(net772),
    .Y(_08626_));
 sky130_fd_sc_hd__and2_2 _09284_ (.A(net474),
    .B(net746),
    .X(_08627_));
 sky130_fd_sc_hd__a22o_2 _09285_ (.A1(net465),
    .A2(net756),
    .B1(net766),
    .B2(net455),
    .X(_08628_));
 sky130_fd_sc_hd__o21ai_4 _09286_ (.A1(_06692_),
    .A2(_08625_),
    .B1(_08628_),
    .Y(_08629_));
 sky130_fd_sc_hd__o2bb2a_2 _09287_ (.A1_N(_08627_),
    .A2_N(_08628_),
    .B1(_06692_),
    .B2(_08625_),
    .X(_08630_));
 sky130_fd_sc_hd__nand2b_2 _09288_ (.A_N(_08630_),
    .B(_08624_),
    .Y(_08631_));
 sky130_fd_sc_hd__xnor2_4 _09289_ (.A(_08624_),
    .B(_08630_),
    .Y(_08632_));
 sky130_fd_sc_hd__nand3_4 _09290_ (.A(_08605_),
    .B(_08612_),
    .C(_08619_),
    .Y(_08633_));
 sky130_fd_sc_hd__nand3_4 _09291_ (.A(_08620_),
    .B(_08632_),
    .C(_08633_),
    .Y(_08634_));
 sky130_fd_sc_hd__nand2_4 _09292_ (.A(_08620_),
    .B(_08634_),
    .Y(_08635_));
 sky130_fd_sc_hd__nor2_1 _09293_ (.A(_06942_),
    .B(_06964_),
    .Y(_08636_));
 sky130_fd_sc_hd__or2_2 _09294_ (.A(_06975_),
    .B(_08636_),
    .X(_08637_));
 sky130_fd_sc_hd__a21o_4 _09295_ (.A1(_08623_),
    .A2(_08631_),
    .B1(_08637_),
    .X(_08638_));
 sky130_fd_sc_hd__nand3_2 _09296_ (.A(_08623_),
    .B(_08631_),
    .C(_08637_),
    .Y(_08639_));
 sky130_fd_sc_hd__o2bb2a_1 _09297_ (.A1_N(net501),
    .A2_N(net711),
    .B1(_06888_),
    .B2(_06899_),
    .X(_08640_));
 sky130_fd_sc_hd__nor2_1 _09298_ (.A(_06909_),
    .B(_08640_),
    .Y(_08641_));
 sky130_fd_sc_hd__and4_1 _09299_ (.A(net481),
    .B(net491),
    .C(net729),
    .D(net737),
    .X(_08642_));
 sky130_fd_sc_hd__a22oi_2 _09300_ (.A1(net492),
    .A2(net730),
    .B1(net737),
    .B2(net482),
    .Y(_08643_));
 sky130_fd_sc_hd__and4bb_1 _09301_ (.A_N(_08642_),
    .B_N(_08643_),
    .C(net501),
    .D(net720),
    .X(_08644_));
 sky130_fd_sc_hd__nor2_1 _09302_ (.A(_08642_),
    .B(_08644_),
    .Y(_08645_));
 sky130_fd_sc_hd__and2b_2 _09303_ (.A_N(_08645_),
    .B(_08641_),
    .X(_08646_));
 sky130_fd_sc_hd__xnor2_1 _09304_ (.A(_08641_),
    .B(_08645_),
    .Y(_08647_));
 sky130_fd_sc_hd__o2bb2a_1 _09305_ (.A1_N(net525),
    .A2_N(net686),
    .B1(_07106_),
    .B2(_07117_),
    .X(_08648_));
 sky130_fd_sc_hd__nor2_1 _09306_ (.A(_07127_),
    .B(_08648_),
    .Y(_08649_));
 sky130_fd_sc_hd__and2_2 _09307_ (.A(_08647_),
    .B(_08649_),
    .X(_08650_));
 sky130_fd_sc_hd__a211o_1 _09308_ (.A1(_08638_),
    .A2(_08639_),
    .B1(_08646_),
    .C1(_08650_),
    .X(_08651_));
 sky130_fd_sc_hd__o211ai_4 _09309_ (.A1(_08646_),
    .A2(_08650_),
    .B1(_08638_),
    .C1(_08639_),
    .Y(_08652_));
 sky130_fd_sc_hd__xnor2_2 _09310_ (.A(_08604_),
    .B(_08635_),
    .Y(_00105_));
 sky130_fd_sc_hd__and3_2 _09311_ (.A(_08651_),
    .B(_08652_),
    .C(_00105_),
    .X(_00106_));
 sky130_fd_sc_hd__a31oi_4 _09312_ (.A1(_06790_),
    .A2(_08603_),
    .A3(_08635_),
    .B1(_00106_),
    .Y(_00107_));
 sky130_fd_sc_hd__or2_2 _09313_ (.A(_08602_),
    .B(_00107_),
    .X(_00108_));
 sky130_fd_sc_hd__xnor2_4 _09314_ (.A(_07269_),
    .B(_07465_),
    .Y(_00109_));
 sky130_fd_sc_hd__a21oi_4 _09315_ (.A1(_08638_),
    .A2(_08652_),
    .B1(_00109_),
    .Y(_00110_));
 sky130_fd_sc_hd__and3_2 _09316_ (.A(_08638_),
    .B(_08652_),
    .C(_00109_),
    .X(_00111_));
 sky130_fd_sc_hd__or3_1 _09317_ (.A(_07182_),
    .B(_07204_),
    .C(_07215_),
    .X(_00112_));
 sky130_fd_sc_hd__nand2_1 _09318_ (.A(_07226_),
    .B(_00112_),
    .Y(_00113_));
 sky130_fd_sc_hd__and4_2 _09319_ (.A(net508),
    .B(net517),
    .C(net703),
    .D(net711),
    .X(_00114_));
 sky130_fd_sc_hd__a22oi_2 _09320_ (.A1(net519),
    .A2(net703),
    .B1(net711),
    .B2(net510),
    .Y(_00115_));
 sky130_fd_sc_hd__and4bb_2 _09321_ (.A_N(_00114_),
    .B_N(_00115_),
    .C(net525),
    .D(net694),
    .X(_00116_));
 sky130_fd_sc_hd__o2bb2a_1 _09322_ (.A1_N(net564),
    .A2_N(net660),
    .B1(_07182_),
    .B2(_07193_),
    .X(_00117_));
 sky130_fd_sc_hd__nor2_2 _09323_ (.A(_07204_),
    .B(_00117_),
    .Y(_00118_));
 sky130_fd_sc_hd__o21ai_4 _09324_ (.A1(_00114_),
    .A2(_00116_),
    .B1(_00118_),
    .Y(_00119_));
 sky130_fd_sc_hd__and4_2 _09325_ (.A(net536),
    .B(net551),
    .C(net679),
    .D(net687),
    .X(_00120_));
 sky130_fd_sc_hd__a22oi_2 _09326_ (.A1(net551),
    .A2(net677),
    .B1(net687),
    .B2(net536),
    .Y(_00121_));
 sky130_fd_sc_hd__and4bb_2 _09327_ (.A_N(_00120_),
    .B_N(_00121_),
    .C(net565),
    .D(net667),
    .X(_00122_));
 sky130_fd_sc_hd__or3_1 _09328_ (.A(_00114_),
    .B(_00116_),
    .C(_00118_),
    .X(_00123_));
 sky130_fd_sc_hd__and2_1 _09329_ (.A(_00119_),
    .B(_00123_),
    .X(_00124_));
 sky130_fd_sc_hd__o21ai_4 _09330_ (.A1(_00120_),
    .A2(_00122_),
    .B1(_00124_),
    .Y(_00125_));
 sky130_fd_sc_hd__a21o_4 _09331_ (.A1(_00119_),
    .A2(_00125_),
    .B1(_00113_),
    .X(_00126_));
 sky130_fd_sc_hd__nand3_2 _09332_ (.A(_00113_),
    .B(_00119_),
    .C(_00125_),
    .Y(_00127_));
 sky130_fd_sc_hd__xnor2_4 _09333_ (.A(_08074_),
    .B(_08085_),
    .Y(_00128_));
 sky130_fd_sc_hd__and3_4 _09334_ (.A(_00126_),
    .B(_00127_),
    .C(_00128_),
    .X(_00129_));
 sky130_fd_sc_hd__inv_2 _09335_ (.A(_00129_),
    .Y(_00130_));
 sky130_fd_sc_hd__o211a_1 _09336_ (.A1(_00110_),
    .A2(_00111_),
    .B1(_00126_),
    .C1(_00130_),
    .X(_00131_));
 sky130_fd_sc_hd__a211oi_4 _09337_ (.A1(_00126_),
    .A2(_00130_),
    .B1(_00110_),
    .C1(_00111_),
    .Y(_00132_));
 sky130_fd_sc_hd__xnor2_2 _09338_ (.A(_08602_),
    .B(_00107_),
    .Y(_00133_));
 sky130_fd_sc_hd__or3_4 _09339_ (.A(_00131_),
    .B(_00132_),
    .C(_00133_),
    .X(_00134_));
 sky130_fd_sc_hd__a21oi_4 _09340_ (.A1(_00108_),
    .A2(_00134_),
    .B1(_08600_),
    .Y(_00135_));
 sky130_fd_sc_hd__a21oi_1 _09341_ (.A1(_08226_),
    .A2(_08247_),
    .B1(_08515_),
    .Y(_00136_));
 sky130_fd_sc_hd__nor2_2 _09342_ (.A(_08521_),
    .B(_00136_),
    .Y(_00137_));
 sky130_fd_sc_hd__o21a_4 _09343_ (.A1(_00110_),
    .A2(_00132_),
    .B1(_00137_),
    .X(_00138_));
 sky130_fd_sc_hd__nor3_4 _09344_ (.A(_00110_),
    .B(_00132_),
    .C(_00137_),
    .Y(_00139_));
 sky130_fd_sc_hd__nor2_1 _09345_ (.A(_08182_),
    .B(_08204_),
    .Y(_00140_));
 sky130_fd_sc_hd__or2_2 _09346_ (.A(_08215_),
    .B(_00140_),
    .X(_00141_));
 sky130_fd_sc_hd__a22oi_4 _09347_ (.A1(net595),
    .A2(\cla_inst.in1[28] ),
    .B1(_08009_),
    .B2(_08020_),
    .Y(_00142_));
 sky130_fd_sc_hd__nor2_2 _09348_ (.A(_08031_),
    .B(_00142_),
    .Y(_00143_));
 sky130_fd_sc_hd__and2_2 _09349_ (.A(net606),
    .B(net661),
    .X(_00144_));
 sky130_fd_sc_hd__and3_2 _09350_ (.A(net581),
    .B(net643),
    .C(_00144_),
    .X(_00145_));
 sky130_fd_sc_hd__a21oi_1 _09351_ (.A1(net581),
    .A2(net661),
    .B1(_07302_),
    .Y(_00146_));
 sky130_fd_sc_hd__and4bb_2 _09352_ (.A_N(_00145_),
    .B_N(_00146_),
    .C(net594),
    .D(net653),
    .X(_00147_));
 sky130_fd_sc_hd__nor2_4 _09353_ (.A(_00145_),
    .B(_00147_),
    .Y(_00148_));
 sky130_fd_sc_hd__or3_4 _09354_ (.A(_08031_),
    .B(_00142_),
    .C(_00148_),
    .X(_00149_));
 sky130_fd_sc_hd__xnor2_4 _09355_ (.A(_00143_),
    .B(_00148_),
    .Y(_00150_));
 sky130_fd_sc_hd__nand2b_1 _09356_ (.A_N(_07596_),
    .B(_00150_),
    .Y(_00151_));
 sky130_fd_sc_hd__nor3_1 _09357_ (.A(_08139_),
    .B(_08161_),
    .C(_08172_),
    .Y(_00152_));
 sky130_fd_sc_hd__or2_1 _09358_ (.A(_08182_),
    .B(_00152_),
    .X(_00153_));
 sky130_fd_sc_hd__a21o_1 _09359_ (.A1(_00149_),
    .A2(_00151_),
    .B1(_00153_),
    .X(_00154_));
 sky130_fd_sc_hd__and3_2 _09360_ (.A(net341),
    .B(net910),
    .C(_08128_),
    .X(_00155_));
 sky130_fd_sc_hd__a21oi_1 _09361_ (.A1(net341),
    .A2(net910),
    .B1(_08128_),
    .Y(_00156_));
 sky130_fd_sc_hd__and4bb_2 _09362_ (.A_N(_00155_),
    .B_N(_00156_),
    .C(net358),
    .D(net892),
    .X(_00157_));
 sky130_fd_sc_hd__o2bb2a_1 _09363_ (.A1_N(net358),
    .A2_N(net881),
    .B1(_08139_),
    .B2(_08150_),
    .X(_00158_));
 sky130_fd_sc_hd__nor2_1 _09364_ (.A(_08161_),
    .B(_00158_),
    .Y(_00159_));
 sky130_fd_sc_hd__o21a_4 _09365_ (.A1(_00155_),
    .A2(_00157_),
    .B1(_00159_),
    .X(_00160_));
 sky130_fd_sc_hd__nand3_1 _09366_ (.A(_00149_),
    .B(_00151_),
    .C(_00153_),
    .Y(_00161_));
 sky130_fd_sc_hd__and2_2 _09367_ (.A(_00154_),
    .B(_00161_),
    .X(_00162_));
 sky130_fd_sc_hd__nand2_1 _09368_ (.A(_00160_),
    .B(_00162_),
    .Y(_00163_));
 sky130_fd_sc_hd__a21o_4 _09369_ (.A1(_00154_),
    .A2(_00163_),
    .B1(_00141_),
    .X(_00164_));
 sky130_fd_sc_hd__nand3_2 _09370_ (.A(_00141_),
    .B(_00154_),
    .C(_00163_),
    .Y(_00165_));
 sky130_fd_sc_hd__nand2_2 _09371_ (.A(net396),
    .B(net811),
    .Y(_00166_));
 sky130_fd_sc_hd__a21oi_2 _09372_ (.A1(net388),
    .A2(net821),
    .B1(_08485_),
    .Y(_00167_));
 sky130_fd_sc_hd__nor2_4 _09373_ (.A(_08491_),
    .B(_00167_),
    .Y(_00168_));
 sky130_fd_sc_hd__o2bb2a_1 _09374_ (.A1_N(net383),
    .A2_N(net842),
    .B1(_08446_),
    .B2(_08454_),
    .X(_00169_));
 sky130_fd_sc_hd__nor2_1 _09375_ (.A(_08461_),
    .B(_00169_),
    .Y(_00170_));
 sky130_fd_sc_hd__and4_1 _09376_ (.A(net371),
    .B(net374),
    .C(net861),
    .D(net871),
    .X(_00171_));
 sky130_fd_sc_hd__a22oi_2 _09377_ (.A1(net380),
    .A2(net861),
    .B1(net871),
    .B2(net371),
    .Y(_00172_));
 sky130_fd_sc_hd__and4bb_1 _09378_ (.A_N(_00171_),
    .B_N(_00172_),
    .C(net381),
    .D(net850),
    .X(_00173_));
 sky130_fd_sc_hd__nor2_1 _09379_ (.A(_00171_),
    .B(_00173_),
    .Y(_00174_));
 sky130_fd_sc_hd__and2b_1 _09380_ (.A_N(_00174_),
    .B(_00170_),
    .X(_00175_));
 sky130_fd_sc_hd__xnor2_1 _09381_ (.A(_00170_),
    .B(_00174_),
    .Y(_00176_));
 sky130_fd_sc_hd__and3_2 _09382_ (.A(net389),
    .B(net830),
    .C(_00176_),
    .X(_00177_));
 sky130_fd_sc_hd__nor2_4 _09383_ (.A(_00175_),
    .B(_00177_),
    .Y(_00178_));
 sky130_fd_sc_hd__and2b_1 _09384_ (.A_N(_00178_),
    .B(_00168_),
    .X(_00179_));
 sky130_fd_sc_hd__xnor2_4 _09385_ (.A(_00168_),
    .B(_00178_),
    .Y(_00180_));
 sky130_fd_sc_hd__xnor2_4 _09386_ (.A(_00166_),
    .B(_00180_),
    .Y(_00181_));
 sky130_fd_sc_hd__and3_4 _09387_ (.A(_00164_),
    .B(_00165_),
    .C(_00181_),
    .X(_00182_));
 sky130_fd_sc_hd__clkinv_2 _09388_ (.A(_00182_),
    .Y(_00183_));
 sky130_fd_sc_hd__a211oi_4 _09389_ (.A1(_00164_),
    .A2(_00183_),
    .B1(_00138_),
    .C1(_00139_),
    .Y(_00184_));
 sky130_fd_sc_hd__o211a_4 _09390_ (.A1(_00138_),
    .A2(_00139_),
    .B1(_00164_),
    .C1(_00183_),
    .X(_00185_));
 sky130_fd_sc_hd__and3_4 _09391_ (.A(_08600_),
    .B(_00108_),
    .C(_00134_),
    .X(_00186_));
 sky130_fd_sc_hd__nor4_4 _09392_ (.A(_00135_),
    .B(net118),
    .C(_00185_),
    .D(_00186_),
    .Y(_00187_));
 sky130_fd_sc_hd__or4_4 _09393_ (.A(_00135_),
    .B(_00184_),
    .C(_00185_),
    .D(_00186_),
    .X(_00188_));
 sky130_fd_sc_hd__o21ai_4 _09394_ (.A1(_00135_),
    .A2(_00187_),
    .B1(_08599_),
    .Y(_00189_));
 sky130_fd_sc_hd__or3_2 _09395_ (.A(_08599_),
    .B(_00135_),
    .C(_00187_),
    .X(_00190_));
 sky130_fd_sc_hd__o211ai_4 _09396_ (.A1(_00138_),
    .A2(net118),
    .B1(_00189_),
    .C1(_00190_),
    .Y(_00191_));
 sky130_fd_sc_hd__a211o_2 _09397_ (.A1(_00189_),
    .A2(_00190_),
    .B1(_00138_),
    .C1(net118),
    .X(_00192_));
 sky130_fd_sc_hd__o22ai_4 _09398_ (.A1(_00184_),
    .A2(_00185_),
    .B1(_00186_),
    .B2(_00135_),
    .Y(_00193_));
 sky130_fd_sc_hd__o21ai_2 _09399_ (.A1(_00131_),
    .A2(_00132_),
    .B1(_00133_),
    .Y(_00194_));
 sky130_fd_sc_hd__a21oi_2 _09400_ (.A1(_08651_),
    .A2(_08652_),
    .B1(_00105_),
    .Y(_00195_));
 sky130_fd_sc_hd__nor2_4 _09401_ (.A(_00106_),
    .B(_00195_),
    .Y(_00196_));
 sky130_fd_sc_hd__a21o_1 _09402_ (.A1(_08620_),
    .A2(_08633_),
    .B1(_08632_),
    .X(_00197_));
 sky130_fd_sc_hd__nand2_2 _09403_ (.A(_08634_),
    .B(_00197_),
    .Y(_00198_));
 sky130_fd_sc_hd__xnor2_2 _09404_ (.A(_08617_),
    .B(_08618_),
    .Y(_00199_));
 sky130_fd_sc_hd__o2bb2a_1 _09405_ (.A1_N(net412),
    .A2_N(net831),
    .B1(_08608_),
    .B2(_08609_),
    .X(_00200_));
 sky130_fd_sc_hd__nor2_2 _09406_ (.A(_08610_),
    .B(_00200_),
    .Y(_00201_));
 sky130_fd_sc_hd__and4_2 _09407_ (.A(net404),
    .B(net419),
    .C(net832),
    .D(net852),
    .X(_00202_));
 sky130_fd_sc_hd__a22oi_2 _09408_ (.A1(net419),
    .A2(net838),
    .B1(net852),
    .B2(net404),
    .Y(_00203_));
 sky130_fd_sc_hd__and4bb_2 _09409_ (.A_N(_00202_),
    .B_N(_00203_),
    .C(net412),
    .D(net841),
    .X(_00204_));
 sky130_fd_sc_hd__nor2_4 _09410_ (.A(_00202_),
    .B(_00204_),
    .Y(_00205_));
 sky130_fd_sc_hd__or3_2 _09411_ (.A(_08610_),
    .B(_00200_),
    .C(_00205_),
    .X(_00206_));
 sky130_fd_sc_hd__nand2_8 _09412_ (.A(net448),
    .B(net793),
    .Y(_00207_));
 sky130_fd_sc_hd__a22oi_4 _09413_ (.A1(net438),
    .A2(net806),
    .B1(net815),
    .B2(net429),
    .Y(_00208_));
 sky130_fd_sc_hd__and4_1 _09414_ (.A(net429),
    .B(net438),
    .C(net801),
    .D(net810),
    .X(_00209_));
 sky130_fd_sc_hd__nor2_2 _09415_ (.A(_00208_),
    .B(_00209_),
    .Y(_00210_));
 sky130_fd_sc_hd__xnor2_4 _09416_ (.A(_00207_),
    .B(_00210_),
    .Y(_00211_));
 sky130_fd_sc_hd__xnor2_4 _09417_ (.A(_00201_),
    .B(_00205_),
    .Y(_00212_));
 sky130_fd_sc_hd__nand2_1 _09418_ (.A(_00211_),
    .B(_00212_),
    .Y(_00213_));
 sky130_fd_sc_hd__a21o_4 _09419_ (.A1(_00206_),
    .A2(_00213_),
    .B1(_00199_),
    .X(_00214_));
 sky130_fd_sc_hd__o21ba_4 _09420_ (.A1(_00207_),
    .A2(_00208_),
    .B1_N(_00209_),
    .X(_00215_));
 sky130_fd_sc_hd__xnor2_4 _09421_ (.A(_08627_),
    .B(_08629_),
    .Y(_00216_));
 sky130_fd_sc_hd__nand2b_2 _09422_ (.A_N(_00215_),
    .B(_00216_),
    .Y(_00217_));
 sky130_fd_sc_hd__xnor2_4 _09423_ (.A(_00215_),
    .B(_00216_),
    .Y(_00218_));
 sky130_fd_sc_hd__and2_4 _09424_ (.A(net472),
    .B(net784),
    .X(_00219_));
 sky130_fd_sc_hd__nand2_8 _09425_ (.A(net465),
    .B(net780),
    .Y(_00220_));
 sky130_fd_sc_hd__nand2_8 _09426_ (.A(net458),
    .B(net782),
    .Y(_00221_));
 sky130_fd_sc_hd__nor2_2 _09427_ (.A(_08626_),
    .B(_00220_),
    .Y(_00222_));
 sky130_fd_sc_hd__nand2_4 _09428_ (.A(net476),
    .B(net758),
    .Y(_00223_));
 sky130_fd_sc_hd__nand2_2 _09429_ (.A(_08625_),
    .B(_00221_),
    .Y(_00224_));
 sky130_fd_sc_hd__and2b_2 _09430_ (.A_N(_00222_),
    .B(_00224_),
    .X(_00225_));
 sky130_fd_sc_hd__a31oi_4 _09431_ (.A1(net476),
    .A2(net759),
    .A3(_00224_),
    .B1(_00222_),
    .Y(_00226_));
 sky130_fd_sc_hd__nand2b_2 _09432_ (.A_N(_00226_),
    .B(_00218_),
    .Y(_00227_));
 sky130_fd_sc_hd__xnor2_4 _09433_ (.A(_00218_),
    .B(_00226_),
    .Y(_00228_));
 sky130_fd_sc_hd__nand3_2 _09434_ (.A(_00199_),
    .B(_00206_),
    .C(_00213_),
    .Y(_00229_));
 sky130_fd_sc_hd__nand3_4 _09435_ (.A(_00214_),
    .B(_00228_),
    .C(_00229_),
    .Y(_00230_));
 sky130_fd_sc_hd__nand2_4 _09436_ (.A(_00214_),
    .B(_00230_),
    .Y(_00231_));
 sky130_fd_sc_hd__and3_2 _09437_ (.A(_08634_),
    .B(_00197_),
    .C(_00231_),
    .X(_00232_));
 sky130_fd_sc_hd__nor2_1 _09438_ (.A(_08647_),
    .B(_08649_),
    .Y(_00233_));
 sky130_fd_sc_hd__or2_2 _09439_ (.A(_08650_),
    .B(_00233_),
    .X(_00234_));
 sky130_fd_sc_hd__a21o_4 _09440_ (.A1(_00217_),
    .A2(_00227_),
    .B1(_00234_),
    .X(_00235_));
 sky130_fd_sc_hd__nand3_2 _09441_ (.A(_00217_),
    .B(_00227_),
    .C(_00234_),
    .Y(_00236_));
 sky130_fd_sc_hd__o2bb2a_1 _09442_ (.A1_N(net501),
    .A2_N(net720),
    .B1(_08642_),
    .B2(_08643_),
    .X(_00237_));
 sky130_fd_sc_hd__nor2_1 _09443_ (.A(_08644_),
    .B(_00237_),
    .Y(_00238_));
 sky130_fd_sc_hd__and4_1 _09444_ (.A(net481),
    .B(net491),
    .C(net737),
    .D(net746),
    .X(_00239_));
 sky130_fd_sc_hd__a22oi_2 _09445_ (.A1(net493),
    .A2(net737),
    .B1(net746),
    .B2(net483),
    .Y(_00240_));
 sky130_fd_sc_hd__and4bb_1 _09446_ (.A_N(_00239_),
    .B_N(_00240_),
    .C(net502),
    .D(net729),
    .X(_00241_));
 sky130_fd_sc_hd__nor2_1 _09447_ (.A(_00239_),
    .B(_00241_),
    .Y(_00242_));
 sky130_fd_sc_hd__and2b_2 _09448_ (.A_N(_00242_),
    .B(_00238_),
    .X(_00243_));
 sky130_fd_sc_hd__xnor2_1 _09449_ (.A(_00238_),
    .B(_00242_),
    .Y(_00244_));
 sky130_fd_sc_hd__o2bb2a_1 _09450_ (.A1_N(net525),
    .A2_N(net695),
    .B1(_00114_),
    .B2(_00115_),
    .X(_00245_));
 sky130_fd_sc_hd__nor2_1 _09451_ (.A(_00116_),
    .B(_00245_),
    .Y(_00246_));
 sky130_fd_sc_hd__and2_2 _09452_ (.A(_00244_),
    .B(_00246_),
    .X(_00247_));
 sky130_fd_sc_hd__a211o_2 _09453_ (.A1(_00235_),
    .A2(_00236_),
    .B1(_00243_),
    .C1(_00247_),
    .X(_00248_));
 sky130_fd_sc_hd__o211ai_4 _09454_ (.A1(_00243_),
    .A2(_00247_),
    .B1(_00235_),
    .C1(_00236_),
    .Y(_00249_));
 sky130_fd_sc_hd__nand2_1 _09455_ (.A(_00248_),
    .B(_00249_),
    .Y(_00250_));
 sky130_fd_sc_hd__xnor2_4 _09456_ (.A(_00198_),
    .B(_00231_),
    .Y(_00251_));
 sky130_fd_sc_hd__a31oi_4 _09457_ (.A1(_00248_),
    .A2(_00249_),
    .A3(_00251_),
    .B1(_00232_),
    .Y(_00252_));
 sky130_fd_sc_hd__and2b_1 _09458_ (.A_N(_00252_),
    .B(_00196_),
    .X(_00253_));
 sky130_fd_sc_hd__a21oi_4 _09459_ (.A1(_00126_),
    .A2(_00127_),
    .B1(_00128_),
    .Y(_00254_));
 sky130_fd_sc_hd__a211o_4 _09460_ (.A1(_00235_),
    .A2(_00249_),
    .B1(_00254_),
    .C1(_00129_),
    .X(_00255_));
 sky130_fd_sc_hd__o211ai_4 _09461_ (.A1(_00129_),
    .A2(_00254_),
    .B1(_00249_),
    .C1(_00235_),
    .Y(_00256_));
 sky130_fd_sc_hd__or3_1 _09462_ (.A(_00120_),
    .B(_00122_),
    .C(_00124_),
    .X(_00257_));
 sky130_fd_sc_hd__nand2_2 _09463_ (.A(_00125_),
    .B(_00257_),
    .Y(_00258_));
 sky130_fd_sc_hd__and4_2 _09464_ (.A(net510),
    .B(net518),
    .C(net714),
    .D(net723),
    .X(_00259_));
 sky130_fd_sc_hd__a22oi_2 _09465_ (.A1(net518),
    .A2(net714),
    .B1(net723),
    .B2(net510),
    .Y(_00260_));
 sky130_fd_sc_hd__and4bb_2 _09466_ (.A_N(_00259_),
    .B_N(_00260_),
    .C(net527),
    .D(net704),
    .X(_00261_));
 sky130_fd_sc_hd__o2bb2a_1 _09467_ (.A1_N(net571),
    .A2_N(net668),
    .B1(_00120_),
    .B2(_00121_),
    .X(_00262_));
 sky130_fd_sc_hd__nor2_2 _09468_ (.A(_00122_),
    .B(_00262_),
    .Y(_00263_));
 sky130_fd_sc_hd__o21ai_4 _09469_ (.A1(_00259_),
    .A2(_00261_),
    .B1(_00263_),
    .Y(_00264_));
 sky130_fd_sc_hd__and4_2 _09470_ (.A(net536),
    .B(net551),
    .C(net687),
    .D(net696),
    .X(_00265_));
 sky130_fd_sc_hd__a22oi_2 _09471_ (.A1(net551),
    .A2(net687),
    .B1(net696),
    .B2(net536),
    .Y(_00266_));
 sky130_fd_sc_hd__and4bb_4 _09472_ (.A_N(_00265_),
    .B_N(_00266_),
    .C(net565),
    .D(net677),
    .X(_00267_));
 sky130_fd_sc_hd__or3_1 _09473_ (.A(_00259_),
    .B(_00261_),
    .C(_00263_),
    .X(_00268_));
 sky130_fd_sc_hd__and2_1 _09474_ (.A(_00264_),
    .B(_00268_),
    .X(_00269_));
 sky130_fd_sc_hd__o21ai_4 _09475_ (.A1(_00265_),
    .A2(_00267_),
    .B1(_00269_),
    .Y(_00270_));
 sky130_fd_sc_hd__a21oi_4 _09476_ (.A1(_00264_),
    .A2(_00270_),
    .B1(_00258_),
    .Y(_00271_));
 sky130_fd_sc_hd__a21o_1 _09477_ (.A1(_00264_),
    .A2(_00270_),
    .B1(_00258_),
    .X(_00272_));
 sky130_fd_sc_hd__nand3_2 _09478_ (.A(_00258_),
    .B(_00264_),
    .C(_00270_),
    .Y(_00273_));
 sky130_fd_sc_hd__xnor2_4 _09479_ (.A(_07596_),
    .B(_00150_),
    .Y(_00274_));
 sky130_fd_sc_hd__and3_4 _09480_ (.A(_00272_),
    .B(_00273_),
    .C(_00274_),
    .X(_00275_));
 sky130_fd_sc_hd__a211o_2 _09481_ (.A1(_00255_),
    .A2(_00256_),
    .B1(_00271_),
    .C1(_00275_),
    .X(_00276_));
 sky130_fd_sc_hd__o211ai_4 _09482_ (.A1(_00271_),
    .A2(_00275_),
    .B1(_00255_),
    .C1(_00256_),
    .Y(_00277_));
 sky130_fd_sc_hd__xnor2_4 _09483_ (.A(_00196_),
    .B(_00252_),
    .Y(_00278_));
 sky130_fd_sc_hd__and3_4 _09484_ (.A(_00276_),
    .B(_00277_),
    .C(_00278_),
    .X(_00279_));
 sky130_fd_sc_hd__o211a_4 _09485_ (.A1(_00253_),
    .A2(_00279_),
    .B1(_00134_),
    .C1(_00194_),
    .X(_00280_));
 sky130_fd_sc_hd__a21oi_4 _09486_ (.A1(_00164_),
    .A2(_00165_),
    .B1(_00181_),
    .Y(_00281_));
 sky130_fd_sc_hd__a211o_4 _09487_ (.A1(_00255_),
    .A2(_00277_),
    .B1(_00281_),
    .C1(_00182_),
    .X(_00282_));
 sky130_fd_sc_hd__o211ai_4 _09488_ (.A1(_00182_),
    .A2(_00281_),
    .B1(_00277_),
    .C1(_00255_),
    .Y(_00283_));
 sky130_fd_sc_hd__xnor2_4 _09489_ (.A(_00160_),
    .B(_00162_),
    .Y(_00284_));
 sky130_fd_sc_hd__o2bb2a_1 _09490_ (.A1_N(net595),
    .A2_N(net653),
    .B1(_00145_),
    .B2(_00146_),
    .X(_00285_));
 sky130_fd_sc_hd__nor2_2 _09491_ (.A(_00147_),
    .B(_00285_),
    .Y(_00286_));
 sky130_fd_sc_hd__and2_2 _09492_ (.A(net607),
    .B(net669),
    .X(_00287_));
 sky130_fd_sc_hd__and3_2 _09493_ (.A(net581),
    .B(net653),
    .C(_00287_),
    .X(_00288_));
 sky130_fd_sc_hd__a21oi_1 _09494_ (.A1(net581),
    .A2(net669),
    .B1(_07987_),
    .Y(_00289_));
 sky130_fd_sc_hd__and4bb_4 _09495_ (.A_N(_00288_),
    .B_N(_00289_),
    .C(net594),
    .D(net661),
    .X(_00290_));
 sky130_fd_sc_hd__o21ai_4 _09496_ (.A1(_00288_),
    .A2(_00290_),
    .B1(_00286_),
    .Y(_00291_));
 sky130_fd_sc_hd__nor3_1 _09497_ (.A(_00155_),
    .B(_00157_),
    .C(_00159_),
    .Y(_00292_));
 sky130_fd_sc_hd__or2_2 _09498_ (.A(_00160_),
    .B(_00292_),
    .X(_00293_));
 sky130_fd_sc_hd__nand2_4 _09499_ (.A(_00291_),
    .B(_00293_),
    .Y(_00294_));
 sky130_fd_sc_hd__or2_4 _09500_ (.A(_00291_),
    .B(_00293_),
    .X(_00295_));
 sky130_fd_sc_hd__nand2_1 _09501_ (.A(net358),
    .B(net911),
    .Y(_00296_));
 sky130_fd_sc_hd__and3_1 _09502_ (.A(net358),
    .B(net910),
    .C(_08128_),
    .X(_00297_));
 sky130_fd_sc_hd__o2bb2a_1 _09503_ (.A1_N(net358),
    .A2_N(net892),
    .B1(_00155_),
    .B2(_00156_),
    .X(_00298_));
 sky130_fd_sc_hd__nor2_1 _09504_ (.A(_00157_),
    .B(_00298_),
    .Y(_00299_));
 sky130_fd_sc_hd__and2_4 _09505_ (.A(_00297_),
    .B(_00299_),
    .X(_00300_));
 sky130_fd_sc_hd__a21boi_4 _09506_ (.A1(_00294_),
    .A2(_00300_),
    .B1_N(_00295_),
    .Y(_00301_));
 sky130_fd_sc_hd__nor2_2 _09507_ (.A(_00284_),
    .B(_00301_),
    .Y(_00302_));
 sky130_fd_sc_hd__xor2_2 _09508_ (.A(_00284_),
    .B(_00301_),
    .X(_00303_));
 sky130_fd_sc_hd__nand2_2 _09509_ (.A(net397),
    .B(net822),
    .Y(_00304_));
 sky130_fd_sc_hd__a21oi_1 _09510_ (.A1(net390),
    .A2(net832),
    .B1(_00176_),
    .Y(_00305_));
 sky130_fd_sc_hd__nor2_1 _09511_ (.A(_00177_),
    .B(_00305_),
    .Y(_00306_));
 sky130_fd_sc_hd__o2bb2a_1 _09512_ (.A1_N(net381),
    .A2_N(net851),
    .B1(_00171_),
    .B2(_00172_),
    .X(_00307_));
 sky130_fd_sc_hd__nor2_1 _09513_ (.A(_00173_),
    .B(_00307_),
    .Y(_00308_));
 sky130_fd_sc_hd__and4_1 _09514_ (.A(net365),
    .B(net374),
    .C(net871),
    .D(net881),
    .X(_00309_));
 sky130_fd_sc_hd__a22oi_2 _09515_ (.A1(net374),
    .A2(net871),
    .B1(net881),
    .B2(net365),
    .Y(_00310_));
 sky130_fd_sc_hd__and4bb_1 _09516_ (.A_N(_00309_),
    .B_N(_00310_),
    .C(net381),
    .D(net861),
    .X(_00311_));
 sky130_fd_sc_hd__nor2_1 _09517_ (.A(_00309_),
    .B(_00311_),
    .Y(_00312_));
 sky130_fd_sc_hd__and2b_1 _09518_ (.A_N(_00312_),
    .B(_00308_),
    .X(_00313_));
 sky130_fd_sc_hd__xnor2_1 _09519_ (.A(_00308_),
    .B(_00312_),
    .Y(_00314_));
 sky130_fd_sc_hd__and3_1 _09520_ (.A(net390),
    .B(net840),
    .C(_00314_),
    .X(_00315_));
 sky130_fd_sc_hd__o21a_1 _09521_ (.A1(_00313_),
    .A2(_00315_),
    .B1(_00306_),
    .X(_00316_));
 sky130_fd_sc_hd__nor3_2 _09522_ (.A(_00306_),
    .B(_00313_),
    .C(_00315_),
    .Y(_00317_));
 sky130_fd_sc_hd__nor2_1 _09523_ (.A(_00316_),
    .B(_00317_),
    .Y(_00318_));
 sky130_fd_sc_hd__xnor2_2 _09524_ (.A(_00304_),
    .B(_00318_),
    .Y(_00319_));
 sky130_fd_sc_hd__and2_2 _09525_ (.A(_00303_),
    .B(_00319_),
    .X(_00320_));
 sky130_fd_sc_hd__o211ai_4 _09526_ (.A1(_00302_),
    .A2(_00320_),
    .B1(_00282_),
    .C1(_00283_),
    .Y(_00321_));
 sky130_fd_sc_hd__a211o_1 _09527_ (.A1(_00282_),
    .A2(_00283_),
    .B1(_00302_),
    .C1(_00320_),
    .X(_00322_));
 sky130_fd_sc_hd__a211oi_1 _09528_ (.A1(_00134_),
    .A2(_00194_),
    .B1(_00253_),
    .C1(_00279_),
    .Y(_00323_));
 sky130_fd_sc_hd__a211o_1 _09529_ (.A1(_00134_),
    .A2(_00194_),
    .B1(_00253_),
    .C1(_00279_),
    .X(_00324_));
 sky130_fd_sc_hd__and4b_4 _09530_ (.A_N(_00280_),
    .B(_00321_),
    .C(_00322_),
    .D(_00324_),
    .X(_00325_));
 sky130_fd_sc_hd__o211a_4 _09531_ (.A1(_00280_),
    .A2(_00325_),
    .B1(_00188_),
    .C1(_00193_),
    .X(_00326_));
 sky130_fd_sc_hd__a211oi_4 _09532_ (.A1(_00188_),
    .A2(_00193_),
    .B1(_00280_),
    .C1(_00325_),
    .Y(_00327_));
 sky130_fd_sc_hd__a211oi_4 _09533_ (.A1(_00282_),
    .A2(_00321_),
    .B1(_00326_),
    .C1(_00327_),
    .Y(_00328_));
 sky130_fd_sc_hd__o211a_2 _09534_ (.A1(_00326_),
    .A2(_00328_),
    .B1(_00191_),
    .C1(_00192_),
    .X(_00329_));
 sky130_fd_sc_hd__a211oi_4 _09535_ (.A1(_00191_),
    .A2(_00192_),
    .B1(_00326_),
    .C1(_00328_),
    .Y(_00330_));
 sky130_fd_sc_hd__nor2_4 _09536_ (.A(_00329_),
    .B(_00330_),
    .Y(_00331_));
 sky130_fd_sc_hd__a31o_4 _09537_ (.A1(net396),
    .A2(net801),
    .A3(_08509_),
    .B1(_08497_),
    .X(_00332_));
 sky130_fd_sc_hd__xor2_4 _09538_ (.A(_00331_),
    .B(_00332_),
    .X(_00333_));
 sky130_fd_sc_hd__o211a_1 _09539_ (.A1(_00326_),
    .A2(_00327_),
    .B1(_00282_),
    .C1(_00321_),
    .X(_00334_));
 sky130_fd_sc_hd__nor2_2 _09540_ (.A(_00328_),
    .B(_00334_),
    .Y(_00335_));
 sky130_fd_sc_hd__o2bb2a_2 _09541_ (.A1_N(_00321_),
    .A2_N(_00322_),
    .B1(_00323_),
    .B2(_00280_),
    .X(_00336_));
 sky130_fd_sc_hd__a21oi_4 _09542_ (.A1(_00276_),
    .A2(_00277_),
    .B1(_00278_),
    .Y(_00337_));
 sky130_fd_sc_hd__xnor2_1 _09543_ (.A(_00250_),
    .B(_00251_),
    .Y(_00338_));
 sky130_fd_sc_hd__a21o_1 _09544_ (.A1(_00214_),
    .A2(_00229_),
    .B1(_00228_),
    .X(_00339_));
 sky130_fd_sc_hd__nand2_1 _09545_ (.A(_00230_),
    .B(_00339_),
    .Y(_00340_));
 sky130_fd_sc_hd__xor2_4 _09546_ (.A(_00211_),
    .B(_00212_),
    .X(_00341_));
 sky130_fd_sc_hd__o2bb2a_1 _09547_ (.A1_N(net412),
    .A2_N(net841),
    .B1(_00202_),
    .B2(_00203_),
    .X(_00342_));
 sky130_fd_sc_hd__nor2_2 _09548_ (.A(_00204_),
    .B(_00342_),
    .Y(_00343_));
 sky130_fd_sc_hd__and4_1 _09549_ (.A(net405),
    .B(net420),
    .C(net845),
    .D(net861),
    .X(_00344_));
 sky130_fd_sc_hd__a22oi_2 _09550_ (.A1(net420),
    .A2(net845),
    .B1(net861),
    .B2(net405),
    .Y(_00345_));
 sky130_fd_sc_hd__and4bb_2 _09551_ (.A_N(_00344_),
    .B_N(_00345_),
    .C(net412),
    .D(net855),
    .X(_00346_));
 sky130_fd_sc_hd__nor2_2 _09552_ (.A(_00344_),
    .B(_00346_),
    .Y(_00347_));
 sky130_fd_sc_hd__and2b_2 _09553_ (.A_N(_00347_),
    .B(_00343_),
    .X(_00348_));
 sky130_fd_sc_hd__a22oi_4 _09554_ (.A1(net438),
    .A2(net815),
    .B1(net822),
    .B2(net429),
    .Y(_00349_));
 sky130_fd_sc_hd__and4_1 _09555_ (.A(net429),
    .B(net438),
    .C(net810),
    .D(net822),
    .X(_00350_));
 sky130_fd_sc_hd__nor2_1 _09556_ (.A(_00349_),
    .B(_00350_),
    .Y(_00351_));
 sky130_fd_sc_hd__nand2_2 _09557_ (.A(net446),
    .B(net801),
    .Y(_00352_));
 sky130_fd_sc_hd__xnor2_2 _09558_ (.A(_00351_),
    .B(_00352_),
    .Y(_00353_));
 sky130_fd_sc_hd__xnor2_2 _09559_ (.A(_00343_),
    .B(_00347_),
    .Y(_00354_));
 sky130_fd_sc_hd__and2_1 _09560_ (.A(_00353_),
    .B(_00354_),
    .X(_00355_));
 sky130_fd_sc_hd__o21ai_4 _09561_ (.A1(_00348_),
    .A2(_00355_),
    .B1(_00341_),
    .Y(_00356_));
 sky130_fd_sc_hd__o21ba_4 _09562_ (.A1(_00349_),
    .A2(_00352_),
    .B1_N(_00350_),
    .X(_00357_));
 sky130_fd_sc_hd__xnor2_4 _09563_ (.A(_00223_),
    .B(_00225_),
    .Y(_00358_));
 sky130_fd_sc_hd__nand2b_2 _09564_ (.A_N(_00357_),
    .B(_00358_),
    .Y(_00359_));
 sky130_fd_sc_hd__xnor2_4 _09565_ (.A(_00357_),
    .B(_00358_),
    .Y(_00360_));
 sky130_fd_sc_hd__nand2_8 _09566_ (.A(net455),
    .B(net793),
    .Y(_00361_));
 sky130_fd_sc_hd__nor2_2 _09567_ (.A(_00220_),
    .B(_00361_),
    .Y(_00362_));
 sky130_fd_sc_hd__nand2_8 _09568_ (.A(net476),
    .B(net771),
    .Y(_00363_));
 sky130_fd_sc_hd__nand2_2 _09569_ (.A(_00220_),
    .B(_00361_),
    .Y(_00364_));
 sky130_fd_sc_hd__and2b_2 _09570_ (.A_N(_00362_),
    .B(_00364_),
    .X(_00365_));
 sky130_fd_sc_hd__a31oi_4 _09571_ (.A1(net477),
    .A2(net770),
    .A3(_00364_),
    .B1(_00362_),
    .Y(_00366_));
 sky130_fd_sc_hd__nand2b_2 _09572_ (.A_N(_00366_),
    .B(_00360_),
    .Y(_00367_));
 sky130_fd_sc_hd__xnor2_2 _09573_ (.A(_00360_),
    .B(_00366_),
    .Y(_00368_));
 sky130_fd_sc_hd__or3_2 _09574_ (.A(_00341_),
    .B(_00348_),
    .C(_00355_),
    .X(_00369_));
 sky130_fd_sc_hd__nand3_2 _09575_ (.A(_00356_),
    .B(_00368_),
    .C(_00369_),
    .Y(_00370_));
 sky130_fd_sc_hd__nand2_2 _09576_ (.A(_00356_),
    .B(_00370_),
    .Y(_00371_));
 sky130_fd_sc_hd__and3_1 _09577_ (.A(_00230_),
    .B(_00339_),
    .C(_00371_),
    .X(_00372_));
 sky130_fd_sc_hd__nor2_1 _09578_ (.A(_00244_),
    .B(_00246_),
    .Y(_00373_));
 sky130_fd_sc_hd__or2_2 _09579_ (.A(_00247_),
    .B(_00373_),
    .X(_00374_));
 sky130_fd_sc_hd__a21o_4 _09580_ (.A1(_00359_),
    .A2(_00367_),
    .B1(_00374_),
    .X(_00375_));
 sky130_fd_sc_hd__nand3_2 _09581_ (.A(_00359_),
    .B(_00367_),
    .C(_00374_),
    .Y(_00376_));
 sky130_fd_sc_hd__o2bb2a_1 _09582_ (.A1_N(net502),
    .A2_N(net729),
    .B1(_00239_),
    .B2(_00240_),
    .X(_00377_));
 sky130_fd_sc_hd__nor2_1 _09583_ (.A(_00241_),
    .B(_00377_),
    .Y(_00378_));
 sky130_fd_sc_hd__and4_1 _09584_ (.A(net483),
    .B(net493),
    .C(net749),
    .D(net755),
    .X(_00379_));
 sky130_fd_sc_hd__a22oi_2 _09585_ (.A1(net493),
    .A2(net749),
    .B1(net755),
    .B2(net483),
    .Y(_00380_));
 sky130_fd_sc_hd__and4bb_1 _09586_ (.A_N(_00379_),
    .B_N(_00380_),
    .C(net502),
    .D(net741),
    .X(_00381_));
 sky130_fd_sc_hd__nor2_1 _09587_ (.A(_00379_),
    .B(_00381_),
    .Y(_00382_));
 sky130_fd_sc_hd__and2b_2 _09588_ (.A_N(_00382_),
    .B(_00378_),
    .X(_00383_));
 sky130_fd_sc_hd__xnor2_1 _09589_ (.A(_00378_),
    .B(_00382_),
    .Y(_00384_));
 sky130_fd_sc_hd__o2bb2a_1 _09590_ (.A1_N(net527),
    .A2_N(net704),
    .B1(_00259_),
    .B2(_00260_),
    .X(_00385_));
 sky130_fd_sc_hd__nor2_1 _09591_ (.A(_00261_),
    .B(_00385_),
    .Y(_00386_));
 sky130_fd_sc_hd__and2_2 _09592_ (.A(_00384_),
    .B(_00386_),
    .X(_00387_));
 sky130_fd_sc_hd__a211o_1 _09593_ (.A1(_00375_),
    .A2(_00376_),
    .B1(_00383_),
    .C1(_00387_),
    .X(_00388_));
 sky130_fd_sc_hd__o211ai_4 _09594_ (.A1(_00383_),
    .A2(_00387_),
    .B1(_00375_),
    .C1(_00376_),
    .Y(_00389_));
 sky130_fd_sc_hd__nand2_1 _09595_ (.A(_00388_),
    .B(_00389_),
    .Y(_00390_));
 sky130_fd_sc_hd__xnor2_2 _09596_ (.A(_00340_),
    .B(_00371_),
    .Y(_00391_));
 sky130_fd_sc_hd__and3_1 _09597_ (.A(_00388_),
    .B(_00389_),
    .C(_00391_),
    .X(_00392_));
 sky130_fd_sc_hd__o21a_1 _09598_ (.A1(_00372_),
    .A2(_00392_),
    .B1(_00338_),
    .X(_00393_));
 sky130_fd_sc_hd__a21oi_4 _09599_ (.A1(_00272_),
    .A2(_00273_),
    .B1(_00274_),
    .Y(_00394_));
 sky130_fd_sc_hd__a211o_4 _09600_ (.A1(_00375_),
    .A2(_00389_),
    .B1(_00394_),
    .C1(_00275_),
    .X(_00395_));
 sky130_fd_sc_hd__o211ai_4 _09601_ (.A1(_00275_),
    .A2(_00394_),
    .B1(_00389_),
    .C1(_00375_),
    .Y(_00396_));
 sky130_fd_sc_hd__or3_1 _09602_ (.A(_00265_),
    .B(_00267_),
    .C(_00269_),
    .X(_00397_));
 sky130_fd_sc_hd__nand2_2 _09603_ (.A(_00270_),
    .B(_00397_),
    .Y(_00398_));
 sky130_fd_sc_hd__and4_1 _09604_ (.A(net510),
    .B(net518),
    .C(net723),
    .D(net732),
    .X(_00399_));
 sky130_fd_sc_hd__a22oi_2 _09605_ (.A1(net518),
    .A2(net723),
    .B1(net732),
    .B2(net510),
    .Y(_00400_));
 sky130_fd_sc_hd__and4bb_1 _09606_ (.A_N(_00399_),
    .B_N(_00400_),
    .C(net527),
    .D(net714),
    .X(_00401_));
 sky130_fd_sc_hd__nor2_2 _09607_ (.A(_00399_),
    .B(_00401_),
    .Y(_00402_));
 sky130_fd_sc_hd__o2bb2a_1 _09608_ (.A1_N(net565),
    .A2_N(net677),
    .B1(_00265_),
    .B2(_00266_),
    .X(_00403_));
 sky130_fd_sc_hd__nor2_1 _09609_ (.A(_00267_),
    .B(_00403_),
    .Y(_00404_));
 sky130_fd_sc_hd__or3_4 _09610_ (.A(_00267_),
    .B(_00402_),
    .C(_00403_),
    .X(_00405_));
 sky130_fd_sc_hd__and4_2 _09611_ (.A(net536),
    .B(net551),
    .C(net696),
    .D(net704),
    .X(_00406_));
 sky130_fd_sc_hd__a22oi_2 _09612_ (.A1(net551),
    .A2(net696),
    .B1(net704),
    .B2(net536),
    .Y(_00407_));
 sky130_fd_sc_hd__and4bb_4 _09613_ (.A_N(_00406_),
    .B_N(_00407_),
    .C(net565),
    .D(net687),
    .X(_00408_));
 sky130_fd_sc_hd__xnor2_2 _09614_ (.A(_00402_),
    .B(_00404_),
    .Y(_00409_));
 sky130_fd_sc_hd__o21ai_4 _09615_ (.A1(_00406_),
    .A2(_00408_),
    .B1(_00409_),
    .Y(_00410_));
 sky130_fd_sc_hd__a21oi_4 _09616_ (.A1(_00405_),
    .A2(_00410_),
    .B1(_00398_),
    .Y(_00411_));
 sky130_fd_sc_hd__a21o_1 _09617_ (.A1(_00405_),
    .A2(_00410_),
    .B1(_00398_),
    .X(_00412_));
 sky130_fd_sc_hd__nand3_2 _09618_ (.A(_00398_),
    .B(_00405_),
    .C(_00410_),
    .Y(_00413_));
 sky130_fd_sc_hd__or3_1 _09619_ (.A(_00286_),
    .B(_00288_),
    .C(_00290_),
    .X(_00414_));
 sky130_fd_sc_hd__and2_2 _09620_ (.A(_00291_),
    .B(_00414_),
    .X(_00415_));
 sky130_fd_sc_hd__and3_4 _09621_ (.A(_00412_),
    .B(_00413_),
    .C(_00415_),
    .X(_00416_));
 sky130_fd_sc_hd__a211o_1 _09622_ (.A1(_00395_),
    .A2(_00396_),
    .B1(_00411_),
    .C1(_00416_),
    .X(_00417_));
 sky130_fd_sc_hd__o211ai_4 _09623_ (.A1(_00411_),
    .A2(_00416_),
    .B1(_00395_),
    .C1(_00396_),
    .Y(_00418_));
 sky130_fd_sc_hd__nor3_1 _09624_ (.A(_00338_),
    .B(_00372_),
    .C(_00392_),
    .Y(_00419_));
 sky130_fd_sc_hd__nor2_1 _09625_ (.A(_00393_),
    .B(_00419_),
    .Y(_00420_));
 sky130_fd_sc_hd__and3_1 _09626_ (.A(_00417_),
    .B(_00418_),
    .C(_00420_),
    .X(_00421_));
 sky130_fd_sc_hd__nor2_2 _09627_ (.A(_00393_),
    .B(_00421_),
    .Y(_00422_));
 sky130_fd_sc_hd__or3_4 _09628_ (.A(_00279_),
    .B(_00337_),
    .C(_00422_),
    .X(_00423_));
 sky130_fd_sc_hd__nand2_2 _09629_ (.A(_00395_),
    .B(_00418_),
    .Y(_00424_));
 sky130_fd_sc_hd__xnor2_1 _09630_ (.A(_00303_),
    .B(_00319_),
    .Y(_00425_));
 sky130_fd_sc_hd__nand2b_2 _09631_ (.A_N(_00425_),
    .B(_00424_),
    .Y(_00426_));
 sky130_fd_sc_hd__xnor2_1 _09632_ (.A(_00424_),
    .B(_00425_),
    .Y(_00427_));
 sky130_fd_sc_hd__a21oi_1 _09633_ (.A1(net390),
    .A2(net842),
    .B1(_00314_),
    .Y(_00428_));
 sky130_fd_sc_hd__nor2_1 _09634_ (.A(_00315_),
    .B(_00428_),
    .Y(_00429_));
 sky130_fd_sc_hd__o2bb2a_1 _09635_ (.A1_N(net381),
    .A2_N(net861),
    .B1(_00309_),
    .B2(_00310_),
    .X(_00430_));
 sky130_fd_sc_hd__nor2_1 _09636_ (.A(_00311_),
    .B(_00430_),
    .Y(_00431_));
 sky130_fd_sc_hd__and4_1 _09637_ (.A(net365),
    .B(net374),
    .C(net881),
    .D(net893),
    .X(_00432_));
 sky130_fd_sc_hd__a22oi_2 _09638_ (.A1(net374),
    .A2(net881),
    .B1(net893),
    .B2(net365),
    .Y(_00433_));
 sky130_fd_sc_hd__and4bb_1 _09639_ (.A_N(_00432_),
    .B_N(_00433_),
    .C(net381),
    .D(net871),
    .X(_00434_));
 sky130_fd_sc_hd__nor2_1 _09640_ (.A(_00432_),
    .B(_00434_),
    .Y(_00435_));
 sky130_fd_sc_hd__and2b_1 _09641_ (.A_N(_00435_),
    .B(_00431_),
    .X(_00436_));
 sky130_fd_sc_hd__xnor2_1 _09642_ (.A(_00431_),
    .B(_00435_),
    .Y(_00437_));
 sky130_fd_sc_hd__and3_1 _09643_ (.A(net390),
    .B(net851),
    .C(_00437_),
    .X(_00438_));
 sky130_fd_sc_hd__o21a_1 _09644_ (.A1(_00436_),
    .A2(_00438_),
    .B1(_00429_),
    .X(_00439_));
 sky130_fd_sc_hd__nor3_1 _09645_ (.A(_00429_),
    .B(_00436_),
    .C(_00438_),
    .Y(_00440_));
 sky130_fd_sc_hd__nor2_1 _09646_ (.A(_00439_),
    .B(_00440_),
    .Y(_00441_));
 sky130_fd_sc_hd__and3_2 _09647_ (.A(net397),
    .B(net832),
    .C(_00441_),
    .X(_00442_));
 sky130_fd_sc_hd__a21oi_2 _09648_ (.A1(net397),
    .A2(net832),
    .B1(_00441_),
    .Y(_00443_));
 sky130_fd_sc_hd__nor2_4 _09649_ (.A(_00442_),
    .B(_00443_),
    .Y(_00444_));
 sky130_fd_sc_hd__o2bb2a_1 _09650_ (.A1_N(net594),
    .A2_N(net661),
    .B1(_00288_),
    .B2(_00289_),
    .X(_00445_));
 sky130_fd_sc_hd__and2_2 _09651_ (.A(net609),
    .B(net677),
    .X(_00446_));
 sky130_fd_sc_hd__and3_1 _09652_ (.A(net581),
    .B(net661),
    .C(_00446_),
    .X(_00447_));
 sky130_fd_sc_hd__a21oi_1 _09653_ (.A1(net581),
    .A2(net677),
    .B1(_00144_),
    .Y(_00448_));
 sky130_fd_sc_hd__and4bb_1 _09654_ (.A_N(_00447_),
    .B_N(_00448_),
    .C(net594),
    .D(net669),
    .X(_00449_));
 sky130_fd_sc_hd__nor2_1 _09655_ (.A(_00447_),
    .B(_00449_),
    .Y(_00450_));
 sky130_fd_sc_hd__or3_4 _09656_ (.A(_00290_),
    .B(_00445_),
    .C(_00450_),
    .X(_00451_));
 sky130_fd_sc_hd__nor2_1 _09657_ (.A(_00297_),
    .B(_00299_),
    .Y(_00452_));
 sky130_fd_sc_hd__or2_2 _09658_ (.A(_00300_),
    .B(_00452_),
    .X(_00453_));
 sky130_fd_sc_hd__nor2_4 _09659_ (.A(_00451_),
    .B(_00453_),
    .Y(_00454_));
 sky130_fd_sc_hd__a211oi_4 _09660_ (.A1(_00294_),
    .A2(_00295_),
    .B1(_00300_),
    .C1(_00454_),
    .Y(_00455_));
 sky130_fd_sc_hd__o211a_1 _09661_ (.A1(_00300_),
    .A2(_00454_),
    .B1(_00294_),
    .C1(_00295_),
    .X(_00456_));
 sky130_fd_sc_hd__nor2_4 _09662_ (.A(_00455_),
    .B(_00456_),
    .Y(_00457_));
 sky130_fd_sc_hd__a32o_1 _09663_ (.A1(_00294_),
    .A2(_00295_),
    .A3(_00454_),
    .B1(_00457_),
    .B2(_00444_),
    .X(_00458_));
 sky130_fd_sc_hd__or2_1 _09664_ (.A(_00427_),
    .B(_00458_),
    .X(_00459_));
 sky130_fd_sc_hd__nand2_2 _09665_ (.A(_00427_),
    .B(_00458_),
    .Y(_00460_));
 sky130_fd_sc_hd__and2_2 _09666_ (.A(_00459_),
    .B(_00460_),
    .X(_00461_));
 sky130_fd_sc_hd__o21ai_4 _09667_ (.A1(_00279_),
    .A2(_00337_),
    .B1(_00422_),
    .Y(_00462_));
 sky130_fd_sc_hd__nand3_4 _09668_ (.A(_00423_),
    .B(_00461_),
    .C(_00462_),
    .Y(_00463_));
 sky130_fd_sc_hd__a211oi_4 _09669_ (.A1(_00423_),
    .A2(_00463_),
    .B1(_00325_),
    .C1(_00336_),
    .Y(_00464_));
 sky130_fd_sc_hd__o211a_2 _09670_ (.A1(_00325_),
    .A2(_00336_),
    .B1(_00423_),
    .C1(_00463_),
    .X(_00465_));
 sky130_fd_sc_hd__a211oi_4 _09671_ (.A1(_00426_),
    .A2(_00460_),
    .B1(_00464_),
    .C1(_00465_),
    .Y(_00466_));
 sky130_fd_sc_hd__o21a_4 _09672_ (.A1(_00464_),
    .A2(_00466_),
    .B1(_00335_),
    .X(_00467_));
 sky130_fd_sc_hd__a31oi_4 _09673_ (.A1(net396),
    .A2(net811),
    .A3(_00180_),
    .B1(_00179_),
    .Y(_00468_));
 sky130_fd_sc_hd__nor3_2 _09674_ (.A(_00335_),
    .B(_00464_),
    .C(_00466_),
    .Y(_00469_));
 sky130_fd_sc_hd__nor3_4 _09675_ (.A(_00467_),
    .B(_00468_),
    .C(_00469_),
    .Y(_00470_));
 sky130_fd_sc_hd__o21ai_2 _09676_ (.A1(_00467_),
    .A2(_00470_),
    .B1(_00333_),
    .Y(_00471_));
 sky130_fd_sc_hd__clkinv_2 _09677_ (.A(_00471_),
    .Y(_00472_));
 sky130_fd_sc_hd__nor3_4 _09678_ (.A(_00333_),
    .B(_00467_),
    .C(_00470_),
    .Y(_00473_));
 sky130_fd_sc_hd__nor2_2 _09679_ (.A(_00472_),
    .B(_00473_),
    .Y(_00474_));
 sky130_fd_sc_hd__o21a_1 _09680_ (.A1(_00467_),
    .A2(_00469_),
    .B1(_00468_),
    .X(_00475_));
 sky130_fd_sc_hd__or2_4 _09681_ (.A(_00470_),
    .B(_00475_),
    .X(_00476_));
 sky130_fd_sc_hd__o211a_1 _09682_ (.A1(_00464_),
    .A2(_00465_),
    .B1(_00426_),
    .C1(_00460_),
    .X(_00477_));
 sky130_fd_sc_hd__a21o_1 _09683_ (.A1(_00423_),
    .A2(_00462_),
    .B1(_00461_),
    .X(_00478_));
 sky130_fd_sc_hd__a21oi_1 _09684_ (.A1(_00417_),
    .A2(_00418_),
    .B1(_00420_),
    .Y(_00479_));
 sky130_fd_sc_hd__nor2_1 _09685_ (.A(_00421_),
    .B(_00479_),
    .Y(_00480_));
 sky130_fd_sc_hd__xnor2_1 _09686_ (.A(_00390_),
    .B(_00391_),
    .Y(_00481_));
 sky130_fd_sc_hd__a21o_1 _09687_ (.A1(_00356_),
    .A2(_00369_),
    .B1(_00368_),
    .X(_00482_));
 sky130_fd_sc_hd__nand2_1 _09688_ (.A(_00370_),
    .B(_00482_),
    .Y(_00483_));
 sky130_fd_sc_hd__xnor2_2 _09689_ (.A(_00353_),
    .B(_00354_),
    .Y(_00484_));
 sky130_fd_sc_hd__o2bb2a_1 _09690_ (.A1_N(net412),
    .A2_N(net852),
    .B1(_00344_),
    .B2(_00345_),
    .X(_00485_));
 sky130_fd_sc_hd__nor2_1 _09691_ (.A(_00346_),
    .B(_00485_),
    .Y(_00486_));
 sky130_fd_sc_hd__and4_1 _09692_ (.A(net405),
    .B(net419),
    .C(net854),
    .D(net871),
    .X(_00487_));
 sky130_fd_sc_hd__a22oi_2 _09693_ (.A1(net421),
    .A2(net854),
    .B1(net874),
    .B2(net405),
    .Y(_00488_));
 sky130_fd_sc_hd__and4bb_2 _09694_ (.A_N(_00487_),
    .B_N(_00488_),
    .C(net418),
    .D(net863),
    .X(_00489_));
 sky130_fd_sc_hd__nor2_2 _09695_ (.A(_00487_),
    .B(_00489_),
    .Y(_00490_));
 sky130_fd_sc_hd__or3_1 _09696_ (.A(_00346_),
    .B(_00485_),
    .C(_00490_),
    .X(_00491_));
 sky130_fd_sc_hd__a22oi_1 _09697_ (.A1(net438),
    .A2(net829),
    .B1(net838),
    .B2(net429),
    .Y(_00492_));
 sky130_fd_sc_hd__and4_2 _09698_ (.A(net429),
    .B(net438),
    .C(net829),
    .D(net838),
    .X(_00493_));
 sky130_fd_sc_hd__nor2_1 _09699_ (.A(_00492_),
    .B(_00493_),
    .Y(_00494_));
 sky130_fd_sc_hd__a21oi_1 _09700_ (.A1(net446),
    .A2(net815),
    .B1(_00494_),
    .Y(_00495_));
 sky130_fd_sc_hd__and3_2 _09701_ (.A(net449),
    .B(net815),
    .C(_00494_),
    .X(_00496_));
 sky130_fd_sc_hd__nor2_2 _09702_ (.A(_00495_),
    .B(_00496_),
    .Y(_00497_));
 sky130_fd_sc_hd__xnor2_2 _09703_ (.A(_00486_),
    .B(_00490_),
    .Y(_00498_));
 sky130_fd_sc_hd__nand2_1 _09704_ (.A(_00497_),
    .B(_00498_),
    .Y(_00499_));
 sky130_fd_sc_hd__a21o_2 _09705_ (.A1(_00491_),
    .A2(_00499_),
    .B1(_00484_),
    .X(_00500_));
 sky130_fd_sc_hd__nor2_4 _09706_ (.A(_00493_),
    .B(_00496_),
    .Y(_00501_));
 sky130_fd_sc_hd__xnor2_4 _09707_ (.A(_00363_),
    .B(_00365_),
    .Y(_00502_));
 sky130_fd_sc_hd__nand2b_2 _09708_ (.A_N(_00501_),
    .B(_00502_),
    .Y(_00503_));
 sky130_fd_sc_hd__xnor2_4 _09709_ (.A(_00501_),
    .B(_00502_),
    .Y(_00504_));
 sky130_fd_sc_hd__nand2_1 _09710_ (.A(net468),
    .B(net806),
    .Y(_00505_));
 sky130_fd_sc_hd__and2_1 _09711_ (.A(net477),
    .B(net780),
    .X(_00506_));
 sky130_fd_sc_hd__nand2_4 _09712_ (.A(net476),
    .B(net780),
    .Y(_00507_));
 sky130_fd_sc_hd__a22o_1 _09713_ (.A1(net465),
    .A2(net793),
    .B1(net806),
    .B2(net455),
    .X(_00508_));
 sky130_fd_sc_hd__o21a_2 _09714_ (.A1(_00361_),
    .A2(_00505_),
    .B1(_00508_),
    .X(_00509_));
 sky130_fd_sc_hd__o2bb2a_2 _09715_ (.A1_N(_00506_),
    .A2_N(_00508_),
    .B1(_00361_),
    .B2(_00505_),
    .X(_00510_));
 sky130_fd_sc_hd__nand2b_2 _09716_ (.A_N(_00510_),
    .B(_00504_),
    .Y(_00511_));
 sky130_fd_sc_hd__xnor2_2 _09717_ (.A(_00504_),
    .B(_00510_),
    .Y(_00512_));
 sky130_fd_sc_hd__nand3_2 _09718_ (.A(_00484_),
    .B(_00491_),
    .C(_00499_),
    .Y(_00513_));
 sky130_fd_sc_hd__nand3_2 _09719_ (.A(_00500_),
    .B(_00512_),
    .C(_00513_),
    .Y(_00514_));
 sky130_fd_sc_hd__nand2_2 _09720_ (.A(_00500_),
    .B(_00514_),
    .Y(_00515_));
 sky130_fd_sc_hd__and3_1 _09721_ (.A(_00370_),
    .B(_00482_),
    .C(_00515_),
    .X(_00516_));
 sky130_fd_sc_hd__nor2_1 _09722_ (.A(_00384_),
    .B(_00386_),
    .Y(_00517_));
 sky130_fd_sc_hd__or2_2 _09723_ (.A(_00387_),
    .B(_00517_),
    .X(_00518_));
 sky130_fd_sc_hd__a21o_4 _09724_ (.A1(_00503_),
    .A2(_00511_),
    .B1(_00518_),
    .X(_00519_));
 sky130_fd_sc_hd__nand3_2 _09725_ (.A(_00503_),
    .B(_00511_),
    .C(_00518_),
    .Y(_00520_));
 sky130_fd_sc_hd__o2bb2a_1 _09726_ (.A1_N(net502),
    .A2_N(net741),
    .B1(_00379_),
    .B2(_00380_),
    .X(_00521_));
 sky130_fd_sc_hd__nor2_1 _09727_ (.A(_00381_),
    .B(_00521_),
    .Y(_00522_));
 sky130_fd_sc_hd__and4_1 _09728_ (.A(net483),
    .B(net493),
    .C(net759),
    .D(net770),
    .X(_00523_));
 sky130_fd_sc_hd__a22oi_2 _09729_ (.A1(net493),
    .A2(net759),
    .B1(net770),
    .B2(net483),
    .Y(_00524_));
 sky130_fd_sc_hd__and4bb_1 _09730_ (.A_N(_00523_),
    .B_N(_00524_),
    .C(net502),
    .D(net749),
    .X(_00525_));
 sky130_fd_sc_hd__nor2_1 _09731_ (.A(_00523_),
    .B(_00525_),
    .Y(_00526_));
 sky130_fd_sc_hd__and2b_2 _09732_ (.A_N(_00526_),
    .B(_00522_),
    .X(_00527_));
 sky130_fd_sc_hd__xnor2_1 _09733_ (.A(_00522_),
    .B(_00526_),
    .Y(_00528_));
 sky130_fd_sc_hd__o2bb2a_1 _09734_ (.A1_N(net527),
    .A2_N(net714),
    .B1(_00399_),
    .B2(_00400_),
    .X(_00529_));
 sky130_fd_sc_hd__nor2_1 _09735_ (.A(_00401_),
    .B(_00529_),
    .Y(_00530_));
 sky130_fd_sc_hd__and2_2 _09736_ (.A(_00528_),
    .B(_00530_),
    .X(_00531_));
 sky130_fd_sc_hd__a211o_1 _09737_ (.A1(_00519_),
    .A2(_00520_),
    .B1(_00527_),
    .C1(_00531_),
    .X(_00532_));
 sky130_fd_sc_hd__o211ai_4 _09738_ (.A1(_00527_),
    .A2(_00531_),
    .B1(_00519_),
    .C1(_00520_),
    .Y(_00533_));
 sky130_fd_sc_hd__xnor2_2 _09739_ (.A(_00483_),
    .B(_00515_),
    .Y(_00534_));
 sky130_fd_sc_hd__and3_1 _09740_ (.A(_00532_),
    .B(_00533_),
    .C(_00534_),
    .X(_00535_));
 sky130_fd_sc_hd__o21a_2 _09741_ (.A1(_00516_),
    .A2(_00535_),
    .B1(_00481_),
    .X(_00536_));
 sky130_fd_sc_hd__inv_2 _09742_ (.A(_00536_),
    .Y(_00537_));
 sky130_fd_sc_hd__a21oi_4 _09743_ (.A1(_00412_),
    .A2(_00413_),
    .B1(_00415_),
    .Y(_00538_));
 sky130_fd_sc_hd__a211o_4 _09744_ (.A1(_00519_),
    .A2(_00533_),
    .B1(_00538_),
    .C1(_00416_),
    .X(_00539_));
 sky130_fd_sc_hd__o211ai_4 _09745_ (.A1(_00416_),
    .A2(_00538_),
    .B1(_00533_),
    .C1(_00519_),
    .Y(_00540_));
 sky130_fd_sc_hd__or3_1 _09746_ (.A(_00406_),
    .B(_00408_),
    .C(_00409_),
    .X(_00541_));
 sky130_fd_sc_hd__nand2_2 _09747_ (.A(_00410_),
    .B(_00541_),
    .Y(_00542_));
 sky130_fd_sc_hd__and4_2 _09748_ (.A(net510),
    .B(net518),
    .C(net732),
    .D(net741),
    .X(_00543_));
 sky130_fd_sc_hd__a22oi_2 _09749_ (.A1(net518),
    .A2(net732),
    .B1(net741),
    .B2(net510),
    .Y(_00544_));
 sky130_fd_sc_hd__and4bb_2 _09750_ (.A_N(_00543_),
    .B_N(_00544_),
    .C(net527),
    .D(net723),
    .X(_00545_));
 sky130_fd_sc_hd__nor2_4 _09751_ (.A(_00543_),
    .B(_00545_),
    .Y(_00546_));
 sky130_fd_sc_hd__o2bb2a_1 _09752_ (.A1_N(net565),
    .A2_N(net687),
    .B1(_00406_),
    .B2(_00407_),
    .X(_00547_));
 sky130_fd_sc_hd__nor2_2 _09753_ (.A(_00408_),
    .B(_00547_),
    .Y(_00548_));
 sky130_fd_sc_hd__or3_4 _09754_ (.A(_00408_),
    .B(_00546_),
    .C(_00547_),
    .X(_00549_));
 sky130_fd_sc_hd__and4_2 _09755_ (.A(net543),
    .B(net557),
    .C(net704),
    .D(net713),
    .X(_00550_));
 sky130_fd_sc_hd__a22oi_2 _09756_ (.A1(net557),
    .A2(net704),
    .B1(net713),
    .B2(net543),
    .Y(_00551_));
 sky130_fd_sc_hd__and4bb_2 _09757_ (.A_N(_00550_),
    .B_N(_00551_),
    .C(net574),
    .D(net696),
    .X(_00552_));
 sky130_fd_sc_hd__xnor2_4 _09758_ (.A(_00546_),
    .B(_00548_),
    .Y(_00553_));
 sky130_fd_sc_hd__o21ai_4 _09759_ (.A1(_00550_),
    .A2(_00552_),
    .B1(_00553_),
    .Y(_00554_));
 sky130_fd_sc_hd__a21oi_4 _09760_ (.A1(_00549_),
    .A2(_00554_),
    .B1(_00542_),
    .Y(_00555_));
 sky130_fd_sc_hd__inv_2 _09761_ (.A(_00555_),
    .Y(_00556_));
 sky130_fd_sc_hd__nand3_2 _09762_ (.A(_00542_),
    .B(_00549_),
    .C(_00554_),
    .Y(_00557_));
 sky130_fd_sc_hd__o21ai_1 _09763_ (.A1(_00290_),
    .A2(_00445_),
    .B1(_00450_),
    .Y(_00558_));
 sky130_fd_sc_hd__and2_1 _09764_ (.A(_00451_),
    .B(_00558_),
    .X(_00559_));
 sky130_fd_sc_hd__and3_4 _09765_ (.A(_00556_),
    .B(_00557_),
    .C(_00559_),
    .X(_00560_));
 sky130_fd_sc_hd__a211o_1 _09766_ (.A1(_00539_),
    .A2(_00540_),
    .B1(_00555_),
    .C1(_00560_),
    .X(_00561_));
 sky130_fd_sc_hd__o211ai_4 _09767_ (.A1(_00555_),
    .A2(_00560_),
    .B1(_00539_),
    .C1(_00540_),
    .Y(_00562_));
 sky130_fd_sc_hd__or3_1 _09768_ (.A(_00481_),
    .B(_00516_),
    .C(_00535_),
    .X(_00563_));
 sky130_fd_sc_hd__and4_2 _09769_ (.A(_00537_),
    .B(_00561_),
    .C(_00562_),
    .D(_00563_),
    .X(_00564_));
 sky130_fd_sc_hd__clkinv_2 _09770_ (.A(_00564_),
    .Y(_00565_));
 sky130_fd_sc_hd__nor2_1 _09771_ (.A(_00536_),
    .B(_00564_),
    .Y(_00566_));
 sky130_fd_sc_hd__and2b_1 _09772_ (.A_N(_00566_),
    .B(_00480_),
    .X(_00567_));
 sky130_fd_sc_hd__or3_2 _09773_ (.A(_00421_),
    .B(_00479_),
    .C(_00566_),
    .X(_00568_));
 sky130_fd_sc_hd__xnor2_4 _09774_ (.A(_00444_),
    .B(_00457_),
    .Y(_00569_));
 sky130_fd_sc_hd__a21oi_4 _09775_ (.A1(_00539_),
    .A2(_00562_),
    .B1(_00569_),
    .Y(_00570_));
 sky130_fd_sc_hd__and3_1 _09776_ (.A(_00539_),
    .B(_00562_),
    .C(_00569_),
    .X(_00571_));
 sky130_fd_sc_hd__nor2_4 _09777_ (.A(_00570_),
    .B(_00571_),
    .Y(_00572_));
 sky130_fd_sc_hd__o2bb2a_1 _09778_ (.A1_N(net594),
    .A2_N(net669),
    .B1(_00447_),
    .B2(_00448_),
    .X(_00573_));
 sky130_fd_sc_hd__and2_2 _09779_ (.A(net607),
    .B(net687),
    .X(_00574_));
 sky130_fd_sc_hd__and3_1 _09780_ (.A(net581),
    .B(net669),
    .C(_00574_),
    .X(_00575_));
 sky130_fd_sc_hd__a21oi_1 _09781_ (.A1(net581),
    .A2(net688),
    .B1(_00287_),
    .Y(_00576_));
 sky130_fd_sc_hd__and4bb_1 _09782_ (.A_N(_00575_),
    .B_N(_00576_),
    .C(net594),
    .D(net677),
    .X(_00577_));
 sky130_fd_sc_hd__nor2_1 _09783_ (.A(_00575_),
    .B(_00577_),
    .Y(_00578_));
 sky130_fd_sc_hd__or3_4 _09784_ (.A(_00449_),
    .B(_00573_),
    .C(_00578_),
    .X(_00579_));
 sky130_fd_sc_hd__a22oi_1 _09785_ (.A1(net358),
    .A2(net901),
    .B1(net910),
    .B2(net356),
    .Y(_00580_));
 sky130_fd_sc_hd__or2_1 _09786_ (.A(_00297_),
    .B(_00580_),
    .X(_00581_));
 sky130_fd_sc_hd__or2_4 _09787_ (.A(_00579_),
    .B(_00581_),
    .X(_00582_));
 sky130_fd_sc_hd__and2_2 _09788_ (.A(_00451_),
    .B(_00453_),
    .X(_00583_));
 sky130_fd_sc_hd__nor2_1 _09789_ (.A(_00454_),
    .B(_00583_),
    .Y(_00584_));
 sky130_fd_sc_hd__xnor2_1 _09790_ (.A(_00582_),
    .B(_00584_),
    .Y(_00585_));
 sky130_fd_sc_hd__nand2_1 _09791_ (.A(net397),
    .B(net842),
    .Y(_00586_));
 sky130_fd_sc_hd__a21oi_1 _09792_ (.A1(net390),
    .A2(net851),
    .B1(_00437_),
    .Y(_00587_));
 sky130_fd_sc_hd__nor2_2 _09793_ (.A(_00438_),
    .B(_00587_),
    .Y(_00588_));
 sky130_fd_sc_hd__o2bb2a_1 _09794_ (.A1_N(net381),
    .A2_N(net871),
    .B1(_00432_),
    .B2(_00433_),
    .X(_00589_));
 sky130_fd_sc_hd__nor2_1 _09795_ (.A(_00434_),
    .B(_00589_),
    .Y(_00590_));
 sky130_fd_sc_hd__and2_1 _09796_ (.A(net374),
    .B(net902),
    .X(_00591_));
 sky130_fd_sc_hd__and3_1 _09797_ (.A(net365),
    .B(net893),
    .C(_00591_),
    .X(_00592_));
 sky130_fd_sc_hd__a22oi_2 _09798_ (.A1(net374),
    .A2(net893),
    .B1(net902),
    .B2(net365),
    .Y(_00593_));
 sky130_fd_sc_hd__and4bb_2 _09799_ (.A_N(_00592_),
    .B_N(_00593_),
    .C(net381),
    .D(net881),
    .X(_00594_));
 sky130_fd_sc_hd__o21a_2 _09800_ (.A1(_00592_),
    .A2(_00594_),
    .B1(_00590_),
    .X(_00595_));
 sky130_fd_sc_hd__nor3_1 _09801_ (.A(_00590_),
    .B(_00592_),
    .C(_00594_),
    .Y(_00596_));
 sky130_fd_sc_hd__nor2_1 _09802_ (.A(_00595_),
    .B(_00596_),
    .Y(_00597_));
 sky130_fd_sc_hd__and3_2 _09803_ (.A(net390),
    .B(net861),
    .C(_00597_),
    .X(_00598_));
 sky130_fd_sc_hd__o21ai_4 _09804_ (.A1(_00595_),
    .A2(_00598_),
    .B1(_00588_),
    .Y(_00599_));
 sky130_fd_sc_hd__or3_1 _09805_ (.A(_00588_),
    .B(_00595_),
    .C(_00598_),
    .X(_00600_));
 sky130_fd_sc_hd__and2_1 _09806_ (.A(_00599_),
    .B(_00600_),
    .X(_00601_));
 sky130_fd_sc_hd__nand2b_2 _09807_ (.A_N(_00586_),
    .B(_00601_),
    .Y(_00602_));
 sky130_fd_sc_hd__xnor2_1 _09808_ (.A(_00586_),
    .B(_00601_),
    .Y(_00603_));
 sky130_fd_sc_hd__nand2_1 _09809_ (.A(_00585_),
    .B(_00603_),
    .Y(_00604_));
 sky130_fd_sc_hd__o31ai_4 _09810_ (.A1(_00454_),
    .A2(_00582_),
    .A3(_00583_),
    .B1(_00604_),
    .Y(_00605_));
 sky130_fd_sc_hd__xor2_4 _09811_ (.A(_00572_),
    .B(_00605_),
    .X(_00606_));
 sky130_fd_sc_hd__or3_2 _09812_ (.A(_00480_),
    .B(_00536_),
    .C(_00564_),
    .X(_00607_));
 sky130_fd_sc_hd__and3_2 _09813_ (.A(_00568_),
    .B(_00606_),
    .C(_00607_),
    .X(_00608_));
 sky130_fd_sc_hd__o211a_1 _09814_ (.A1(_00567_),
    .A2(_00608_),
    .B1(_00463_),
    .C1(_00478_),
    .X(_00609_));
 sky130_fd_sc_hd__a21o_2 _09815_ (.A1(_00572_),
    .A2(_00605_),
    .B1(_00570_),
    .X(_00610_));
 sky130_fd_sc_hd__a211o_1 _09816_ (.A1(_00463_),
    .A2(_00478_),
    .B1(_00567_),
    .C1(_00608_),
    .X(_00611_));
 sky130_fd_sc_hd__and2b_1 _09817_ (.A_N(_00609_),
    .B(_00611_),
    .X(_00612_));
 sky130_fd_sc_hd__a21oi_1 _09818_ (.A1(_00610_),
    .A2(_00611_),
    .B1(_00609_),
    .Y(_00613_));
 sky130_fd_sc_hd__nor3_1 _09819_ (.A(_00466_),
    .B(_00477_),
    .C(_00613_),
    .Y(_00614_));
 sky130_fd_sc_hd__o21ba_4 _09820_ (.A1(_00304_),
    .A2(_00317_),
    .B1_N(_00316_),
    .X(_00615_));
 sky130_fd_sc_hd__o21a_1 _09821_ (.A1(_00466_),
    .A2(_00477_),
    .B1(_00613_),
    .X(_00616_));
 sky130_fd_sc_hd__nor2_2 _09822_ (.A(_00614_),
    .B(_00616_),
    .Y(_00617_));
 sky130_fd_sc_hd__o21ba_2 _09823_ (.A1(_00615_),
    .A2(_00616_),
    .B1_N(_00614_),
    .X(_00618_));
 sky130_fd_sc_hd__nor2_4 _09824_ (.A(_00476_),
    .B(_00618_),
    .Y(_00619_));
 sky130_fd_sc_hd__and2_1 _09825_ (.A(_00476_),
    .B(_00618_),
    .X(_00620_));
 sky130_fd_sc_hd__nor2_1 _09826_ (.A(_00619_),
    .B(_00620_),
    .Y(_00621_));
 sky130_fd_sc_hd__xnor2_4 _09827_ (.A(_00615_),
    .B(_00617_),
    .Y(_00622_));
 sky130_fd_sc_hd__xor2_2 _09828_ (.A(_00610_),
    .B(_00612_),
    .X(_00623_));
 sky130_fd_sc_hd__a21oi_4 _09829_ (.A1(_00568_),
    .A2(_00607_),
    .B1(_00606_),
    .Y(_00624_));
 sky130_fd_sc_hd__a22o_2 _09830_ (.A1(_00561_),
    .A2(_00562_),
    .B1(_00563_),
    .B2(_00537_),
    .X(_00625_));
 sky130_fd_sc_hd__a21oi_1 _09831_ (.A1(_00532_),
    .A2(_00533_),
    .B1(_00534_),
    .Y(_00626_));
 sky130_fd_sc_hd__nor2_1 _09832_ (.A(_00535_),
    .B(_00626_),
    .Y(_00627_));
 sky130_fd_sc_hd__a21o_1 _09833_ (.A1(_00500_),
    .A2(_00513_),
    .B1(_00512_),
    .X(_00628_));
 sky130_fd_sc_hd__nand2_2 _09834_ (.A(_00514_),
    .B(_00628_),
    .Y(_00629_));
 sky130_fd_sc_hd__xnor2_2 _09835_ (.A(_00497_),
    .B(_00498_),
    .Y(_00630_));
 sky130_fd_sc_hd__o2bb2a_1 _09836_ (.A1_N(net418),
    .A2_N(net864),
    .B1(_00487_),
    .B2(_00488_),
    .X(_00631_));
 sky130_fd_sc_hd__nor2_2 _09837_ (.A(_00489_),
    .B(_00631_),
    .Y(_00632_));
 sky130_fd_sc_hd__and4_2 _09838_ (.A(net406),
    .B(net422),
    .C(net863),
    .D(net882),
    .X(_00633_));
 sky130_fd_sc_hd__a22oi_2 _09839_ (.A1(net422),
    .A2(net863),
    .B1(net882),
    .B2(net406),
    .Y(_00634_));
 sky130_fd_sc_hd__and4bb_4 _09840_ (.A_N(_00633_),
    .B_N(_00634_),
    .C(net414),
    .D(net872),
    .X(_00635_));
 sky130_fd_sc_hd__nor2_4 _09841_ (.A(_00633_),
    .B(_00635_),
    .Y(_00636_));
 sky130_fd_sc_hd__or3_1 _09842_ (.A(_00489_),
    .B(_00631_),
    .C(_00636_),
    .X(_00637_));
 sky130_fd_sc_hd__and4_1 _09843_ (.A(net435),
    .B(net441),
    .C(net833),
    .D(net843),
    .X(_00638_));
 sky130_fd_sc_hd__a22oi_4 _09844_ (.A1(net441),
    .A2(net833),
    .B1(net843),
    .B2(net435),
    .Y(_00639_));
 sky130_fd_sc_hd__nor2_2 _09845_ (.A(_00638_),
    .B(_00639_),
    .Y(_00640_));
 sky130_fd_sc_hd__nand2_4 _09846_ (.A(net449),
    .B(net826),
    .Y(_00641_));
 sky130_fd_sc_hd__xnor2_4 _09847_ (.A(_00640_),
    .B(_00641_),
    .Y(_00642_));
 sky130_fd_sc_hd__xnor2_4 _09848_ (.A(_00632_),
    .B(_00636_),
    .Y(_00643_));
 sky130_fd_sc_hd__nand2_1 _09849_ (.A(_00642_),
    .B(_00643_),
    .Y(_00644_));
 sky130_fd_sc_hd__a21o_2 _09850_ (.A1(_00637_),
    .A2(_00644_),
    .B1(_00630_),
    .X(_00645_));
 sky130_fd_sc_hd__o21ba_4 _09851_ (.A1(_00639_),
    .A2(_00641_),
    .B1_N(_00638_),
    .X(_00646_));
 sky130_fd_sc_hd__xnor2_4 _09852_ (.A(_00507_),
    .B(_00509_),
    .Y(_00647_));
 sky130_fd_sc_hd__nand2b_1 _09853_ (.A_N(_00646_),
    .B(_00647_),
    .Y(_00648_));
 sky130_fd_sc_hd__xnor2_4 _09854_ (.A(_00646_),
    .B(_00647_),
    .Y(_00649_));
 sky130_fd_sc_hd__and4_1 _09855_ (.A(net458),
    .B(net468),
    .C(net806),
    .D(net815),
    .X(_00650_));
 sky130_fd_sc_hd__nand2_1 _09856_ (.A(net458),
    .B(net815),
    .Y(_00651_));
 sky130_fd_sc_hd__a21o_2 _09857_ (.A1(_00505_),
    .A2(_00651_),
    .B1(_00650_),
    .X(_00652_));
 sky130_fd_sc_hd__and2_4 _09858_ (.A(net477),
    .B(net792),
    .X(_00653_));
 sky130_fd_sc_hd__nand2_8 _09859_ (.A(net478),
    .B(net797),
    .Y(_00654_));
 sky130_fd_sc_hd__o21ba_2 _09860_ (.A1(_00652_),
    .A2(_00654_),
    .B1_N(_00650_),
    .X(_00655_));
 sky130_fd_sc_hd__nand2b_1 _09861_ (.A_N(_00655_),
    .B(_00649_),
    .Y(_00656_));
 sky130_fd_sc_hd__xnor2_2 _09862_ (.A(_00649_),
    .B(_00655_),
    .Y(_00657_));
 sky130_fd_sc_hd__nand3_2 _09863_ (.A(_00630_),
    .B(_00637_),
    .C(_00644_),
    .Y(_00658_));
 sky130_fd_sc_hd__nand3_4 _09864_ (.A(_00645_),
    .B(_00657_),
    .C(_00658_),
    .Y(_00659_));
 sky130_fd_sc_hd__nand2_4 _09865_ (.A(_00645_),
    .B(_00659_),
    .Y(_00660_));
 sky130_fd_sc_hd__and3_1 _09866_ (.A(_00514_),
    .B(_00628_),
    .C(_00660_),
    .X(_00661_));
 sky130_fd_sc_hd__nor2_1 _09867_ (.A(_00528_),
    .B(_00530_),
    .Y(_00662_));
 sky130_fd_sc_hd__or2_2 _09868_ (.A(_00531_),
    .B(_00662_),
    .X(_00663_));
 sky130_fd_sc_hd__a21o_2 _09869_ (.A1(_00648_),
    .A2(_00656_),
    .B1(_00663_),
    .X(_00664_));
 sky130_fd_sc_hd__nand3_2 _09870_ (.A(_00648_),
    .B(_00656_),
    .C(_00663_),
    .Y(_00665_));
 sky130_fd_sc_hd__o2bb2a_1 _09871_ (.A1_N(net502),
    .A2_N(net749),
    .B1(_00523_),
    .B2(_00524_),
    .X(_00666_));
 sky130_fd_sc_hd__nor2_2 _09872_ (.A(_00525_),
    .B(_00666_),
    .Y(_00667_));
 sky130_fd_sc_hd__and4_1 _09873_ (.A(net483),
    .B(net493),
    .C(net770),
    .D(net780),
    .X(_00668_));
 sky130_fd_sc_hd__a22oi_2 _09874_ (.A1(net499),
    .A2(net770),
    .B1(net780),
    .B2(net489),
    .Y(_00669_));
 sky130_fd_sc_hd__and4bb_2 _09875_ (.A_N(_00668_),
    .B_N(_00669_),
    .C(net506),
    .D(net759),
    .X(_00670_));
 sky130_fd_sc_hd__nor2_2 _09876_ (.A(_00668_),
    .B(_00670_),
    .Y(_00671_));
 sky130_fd_sc_hd__and2b_2 _09877_ (.A_N(_00671_),
    .B(_00667_),
    .X(_00672_));
 sky130_fd_sc_hd__xnor2_2 _09878_ (.A(_00667_),
    .B(_00671_),
    .Y(_00673_));
 sky130_fd_sc_hd__o2bb2a_1 _09879_ (.A1_N(net527),
    .A2_N(net723),
    .B1(_00543_),
    .B2(_00544_),
    .X(_00674_));
 sky130_fd_sc_hd__nor2_2 _09880_ (.A(_00545_),
    .B(_00674_),
    .Y(_00675_));
 sky130_fd_sc_hd__and2_2 _09881_ (.A(_00673_),
    .B(_00675_),
    .X(_00676_));
 sky130_fd_sc_hd__o211ai_4 _09882_ (.A1(_00672_),
    .A2(_00676_),
    .B1(_00664_),
    .C1(_00665_),
    .Y(_00677_));
 sky130_fd_sc_hd__a211o_2 _09883_ (.A1(_00664_),
    .A2(_00665_),
    .B1(_00672_),
    .C1(_00676_),
    .X(_00678_));
 sky130_fd_sc_hd__xnor2_4 _09884_ (.A(_00629_),
    .B(_00660_),
    .Y(_00679_));
 sky130_fd_sc_hd__and3_2 _09885_ (.A(_00677_),
    .B(_00678_),
    .C(_00679_),
    .X(_00680_));
 sky130_fd_sc_hd__o21a_2 _09886_ (.A1(_00661_),
    .A2(_00680_),
    .B1(_00627_),
    .X(_00681_));
 sky130_fd_sc_hd__a21oi_2 _09887_ (.A1(_00556_),
    .A2(_00557_),
    .B1(_00559_),
    .Y(_00682_));
 sky130_fd_sc_hd__a211oi_2 _09888_ (.A1(_00664_),
    .A2(_00677_),
    .B1(_00682_),
    .C1(_00560_),
    .Y(_00683_));
 sky130_fd_sc_hd__o211a_1 _09889_ (.A1(_00560_),
    .A2(_00682_),
    .B1(_00677_),
    .C1(_00664_),
    .X(_00684_));
 sky130_fd_sc_hd__or3_1 _09890_ (.A(_00550_),
    .B(_00552_),
    .C(_00553_),
    .X(_00685_));
 sky130_fd_sc_hd__nand2_1 _09891_ (.A(_00554_),
    .B(_00685_),
    .Y(_00686_));
 sky130_fd_sc_hd__and4_1 _09892_ (.A(net514),
    .B(net521),
    .C(net741),
    .D(net749),
    .X(_00687_));
 sky130_fd_sc_hd__a22oi_2 _09893_ (.A1(net521),
    .A2(net741),
    .B1(net749),
    .B2(net514),
    .Y(_00688_));
 sky130_fd_sc_hd__and4bb_2 _09894_ (.A_N(_00687_),
    .B_N(_00688_),
    .C(net531),
    .D(net731),
    .X(_00689_));
 sky130_fd_sc_hd__nor2_2 _09895_ (.A(_00687_),
    .B(_00689_),
    .Y(_00690_));
 sky130_fd_sc_hd__o2bb2a_1 _09896_ (.A1_N(net565),
    .A2_N(net696),
    .B1(_00550_),
    .B2(_00551_),
    .X(_00691_));
 sky130_fd_sc_hd__nor2_1 _09897_ (.A(_00552_),
    .B(_00691_),
    .Y(_00692_));
 sky130_fd_sc_hd__or3_1 _09898_ (.A(_00552_),
    .B(_00690_),
    .C(_00691_),
    .X(_00693_));
 sky130_fd_sc_hd__and4_2 _09899_ (.A(net543),
    .B(net557),
    .C(net713),
    .D(net722),
    .X(_00694_));
 sky130_fd_sc_hd__a22oi_2 _09900_ (.A1(net557),
    .A2(net713),
    .B1(net722),
    .B2(net543),
    .Y(_00695_));
 sky130_fd_sc_hd__and4bb_2 _09901_ (.A_N(_00694_),
    .B_N(_00695_),
    .C(net574),
    .D(net705),
    .X(_00696_));
 sky130_fd_sc_hd__xnor2_2 _09902_ (.A(_00690_),
    .B(_00692_),
    .Y(_00697_));
 sky130_fd_sc_hd__o21ai_2 _09903_ (.A1(_00694_),
    .A2(_00696_),
    .B1(_00697_),
    .Y(_00698_));
 sky130_fd_sc_hd__a21o_1 _09904_ (.A1(_00693_),
    .A2(_00698_),
    .B1(_00686_),
    .X(_00699_));
 sky130_fd_sc_hd__inv_2 _09905_ (.A(_00699_),
    .Y(_00700_));
 sky130_fd_sc_hd__nand3_1 _09906_ (.A(_00686_),
    .B(_00693_),
    .C(_00698_),
    .Y(_00701_));
 sky130_fd_sc_hd__o21ai_1 _09907_ (.A1(_00449_),
    .A2(_00573_),
    .B1(_00578_),
    .Y(_00702_));
 sky130_fd_sc_hd__and2_1 _09908_ (.A(_00579_),
    .B(_00702_),
    .X(_00703_));
 sky130_fd_sc_hd__and3_1 _09909_ (.A(_00699_),
    .B(_00701_),
    .C(_00703_),
    .X(_00704_));
 sky130_fd_sc_hd__nor2_1 _09910_ (.A(_00700_),
    .B(_00704_),
    .Y(_00705_));
 sky130_fd_sc_hd__o21ai_1 _09911_ (.A1(_00683_),
    .A2(_00684_),
    .B1(_00705_),
    .Y(_00706_));
 sky130_fd_sc_hd__or3_1 _09912_ (.A(_00683_),
    .B(_00684_),
    .C(_00705_),
    .X(_00707_));
 sky130_fd_sc_hd__nand2_2 _09913_ (.A(_00706_),
    .B(_00707_),
    .Y(_00708_));
 sky130_fd_sc_hd__nor3_1 _09914_ (.A(_00627_),
    .B(_00661_),
    .C(_00680_),
    .Y(_00709_));
 sky130_fd_sc_hd__or2_2 _09915_ (.A(_00681_),
    .B(_00709_),
    .X(_00710_));
 sky130_fd_sc_hd__nor2_4 _09916_ (.A(_00708_),
    .B(_00710_),
    .Y(_00711_));
 sky130_fd_sc_hd__o211ai_4 _09917_ (.A1(_00681_),
    .A2(_00711_),
    .B1(_00565_),
    .C1(_00625_),
    .Y(_00712_));
 sky130_fd_sc_hd__o21bai_2 _09918_ (.A1(_00684_),
    .A2(_00705_),
    .B1_N(_00683_),
    .Y(_00713_));
 sky130_fd_sc_hd__or2_1 _09919_ (.A(_00585_),
    .B(_00603_),
    .X(_00714_));
 sky130_fd_sc_hd__and2_1 _09920_ (.A(_00604_),
    .B(_00714_),
    .X(_00715_));
 sky130_fd_sc_hd__nand2_2 _09921_ (.A(_00713_),
    .B(_00715_),
    .Y(_00716_));
 sky130_fd_sc_hd__or2_1 _09922_ (.A(_00713_),
    .B(_00715_),
    .X(_00717_));
 sky130_fd_sc_hd__and2_1 _09923_ (.A(_00716_),
    .B(_00717_),
    .X(_00718_));
 sky130_fd_sc_hd__o2bb2a_1 _09924_ (.A1_N(net594),
    .A2_N(net677),
    .B1(_00575_),
    .B2(_00576_),
    .X(_00719_));
 sky130_fd_sc_hd__and2_2 _09925_ (.A(net607),
    .B(net697),
    .X(_00720_));
 sky130_fd_sc_hd__and3_1 _09926_ (.A(net582),
    .B(net677),
    .C(_00720_),
    .X(_00721_));
 sky130_fd_sc_hd__a21oi_1 _09927_ (.A1(net582),
    .A2(net696),
    .B1(_00446_),
    .Y(_00722_));
 sky130_fd_sc_hd__and4bb_1 _09928_ (.A_N(_00721_),
    .B_N(_00722_),
    .C(net595),
    .D(net687),
    .X(_00723_));
 sky130_fd_sc_hd__nor2_1 _09929_ (.A(_00721_),
    .B(_00723_),
    .Y(_00724_));
 sky130_fd_sc_hd__or3_4 _09930_ (.A(_00577_),
    .B(_00719_),
    .C(_00724_),
    .X(_00725_));
 sky130_fd_sc_hd__or2_1 _09931_ (.A(_00296_),
    .B(_00725_),
    .X(_00726_));
 sky130_fd_sc_hd__nand2_1 _09932_ (.A(_00579_),
    .B(_00581_),
    .Y(_00727_));
 sky130_fd_sc_hd__nand2_1 _09933_ (.A(_00582_),
    .B(_00727_),
    .Y(_00728_));
 sky130_fd_sc_hd__nor2_1 _09934_ (.A(_00726_),
    .B(_00728_),
    .Y(_00729_));
 sky130_fd_sc_hd__and2_1 _09935_ (.A(_00726_),
    .B(_00728_),
    .X(_00730_));
 sky130_fd_sc_hd__nor2_2 _09936_ (.A(_00729_),
    .B(_00730_),
    .Y(_00731_));
 sky130_fd_sc_hd__nand2_2 _09937_ (.A(net398),
    .B(net854),
    .Y(_00732_));
 sky130_fd_sc_hd__a21oi_1 _09938_ (.A1(net390),
    .A2(net861),
    .B1(_00597_),
    .Y(_00733_));
 sky130_fd_sc_hd__nor2_1 _09939_ (.A(_00598_),
    .B(_00733_),
    .Y(_00734_));
 sky130_fd_sc_hd__o2bb2a_1 _09940_ (.A1_N(net382),
    .A2_N(net881),
    .B1(_00592_),
    .B2(_00593_),
    .X(_00735_));
 sky130_fd_sc_hd__nor2_2 _09941_ (.A(_00594_),
    .B(_00735_),
    .Y(_00736_));
 sky130_fd_sc_hd__and3_1 _09942_ (.A(net365),
    .B(net911),
    .C(_00591_),
    .X(_00737_));
 sky130_fd_sc_hd__a21oi_1 _09943_ (.A1(net365),
    .A2(net911),
    .B1(_00591_),
    .Y(_00738_));
 sky130_fd_sc_hd__and4bb_1 _09944_ (.A_N(_00737_),
    .B_N(_00738_),
    .C(net381),
    .D(net893),
    .X(_00739_));
 sky130_fd_sc_hd__nor2_2 _09945_ (.A(_00737_),
    .B(_00739_),
    .Y(_00740_));
 sky130_fd_sc_hd__and2b_1 _09946_ (.A_N(_00740_),
    .B(_00736_),
    .X(_00741_));
 sky130_fd_sc_hd__nand2_1 _09947_ (.A(net391),
    .B(net872),
    .Y(_00742_));
 sky130_fd_sc_hd__xnor2_2 _09948_ (.A(_00736_),
    .B(_00740_),
    .Y(_00743_));
 sky130_fd_sc_hd__and3_1 _09949_ (.A(net391),
    .B(net872),
    .C(_00743_),
    .X(_00744_));
 sky130_fd_sc_hd__o21a_2 _09950_ (.A1(_00741_),
    .A2(_00744_),
    .B1(_00734_),
    .X(_00745_));
 sky130_fd_sc_hd__nor3_2 _09951_ (.A(_00734_),
    .B(_00741_),
    .C(_00744_),
    .Y(_00746_));
 sky130_fd_sc_hd__nor2_4 _09952_ (.A(_00745_),
    .B(_00746_),
    .Y(_00747_));
 sky130_fd_sc_hd__xnor2_4 _09953_ (.A(_00732_),
    .B(_00747_),
    .Y(_00748_));
 sky130_fd_sc_hd__a21o_1 _09954_ (.A1(_00731_),
    .A2(_00748_),
    .B1(_00729_),
    .X(_00749_));
 sky130_fd_sc_hd__nand2_2 _09955_ (.A(_00718_),
    .B(_00749_),
    .Y(_00750_));
 sky130_fd_sc_hd__or2_1 _09956_ (.A(_00718_),
    .B(_00749_),
    .X(_00751_));
 sky130_fd_sc_hd__and2_2 _09957_ (.A(_00750_),
    .B(_00751_),
    .X(_00752_));
 sky130_fd_sc_hd__a211o_4 _09958_ (.A1(_00565_),
    .A2(_00625_),
    .B1(_00681_),
    .C1(_00711_),
    .X(_00753_));
 sky130_fd_sc_hd__and3_2 _09959_ (.A(_00712_),
    .B(_00752_),
    .C(_00753_),
    .X(_00754_));
 sky130_fd_sc_hd__nand3_2 _09960_ (.A(_00712_),
    .B(_00752_),
    .C(_00753_),
    .Y(_00755_));
 sky130_fd_sc_hd__a211oi_4 _09961_ (.A1(_00712_),
    .A2(_00755_),
    .B1(_00608_),
    .C1(_00624_),
    .Y(_00756_));
 sky130_fd_sc_hd__o211a_2 _09962_ (.A1(_00608_),
    .A2(_00624_),
    .B1(_00712_),
    .C1(_00755_),
    .X(_00757_));
 sky130_fd_sc_hd__a211oi_4 _09963_ (.A1(_00716_),
    .A2(_00750_),
    .B1(_00756_),
    .C1(_00757_),
    .Y(_00758_));
 sky130_fd_sc_hd__nor2_1 _09964_ (.A(_00756_),
    .B(_00758_),
    .Y(_00759_));
 sky130_fd_sc_hd__and2b_2 _09965_ (.A_N(_00759_),
    .B(_00623_),
    .X(_00760_));
 sky130_fd_sc_hd__xnor2_1 _09966_ (.A(_00623_),
    .B(_00759_),
    .Y(_00761_));
 sky130_fd_sc_hd__o21a_2 _09967_ (.A1(_00439_),
    .A2(_00442_),
    .B1(_00761_),
    .X(_00762_));
 sky130_fd_sc_hd__or3_4 _09968_ (.A(_00622_),
    .B(_00760_),
    .C(_00762_),
    .X(_00763_));
 sky130_fd_sc_hd__nor3_1 _09969_ (.A(_00439_),
    .B(_00442_),
    .C(_00761_),
    .Y(_00764_));
 sky130_fd_sc_hd__or2_2 _09970_ (.A(_00762_),
    .B(_00764_),
    .X(_00765_));
 sky130_fd_sc_hd__o211a_2 _09971_ (.A1(_00756_),
    .A2(_00757_),
    .B1(_00716_),
    .C1(_00750_),
    .X(_00766_));
 sky130_fd_sc_hd__a21oi_4 _09972_ (.A1(_00712_),
    .A2(_00753_),
    .B1(_00752_),
    .Y(_00767_));
 sky130_fd_sc_hd__and2_2 _09973_ (.A(_00708_),
    .B(_00710_),
    .X(_00768_));
 sky130_fd_sc_hd__a21oi_4 _09974_ (.A1(_00677_),
    .A2(_00678_),
    .B1(_00679_),
    .Y(_00769_));
 sky130_fd_sc_hd__a21o_1 _09975_ (.A1(_00645_),
    .A2(_00658_),
    .B1(_00657_),
    .X(_00770_));
 sky130_fd_sc_hd__xnor2_4 _09976_ (.A(_00642_),
    .B(_00643_),
    .Y(_00771_));
 sky130_fd_sc_hd__o2bb2a_1 _09977_ (.A1_N(net414),
    .A2_N(net872),
    .B1(_00633_),
    .B2(_00634_),
    .X(_00772_));
 sky130_fd_sc_hd__nor2_2 _09978_ (.A(_00635_),
    .B(_00772_),
    .Y(_00773_));
 sky130_fd_sc_hd__and4_2 _09979_ (.A(net406),
    .B(net422),
    .C(net872),
    .D(net894),
    .X(_00774_));
 sky130_fd_sc_hd__a22oi_2 _09980_ (.A1(net422),
    .A2(net872),
    .B1(net894),
    .B2(net406),
    .Y(_00775_));
 sky130_fd_sc_hd__and4bb_4 _09981_ (.A_N(_00774_),
    .B_N(_00775_),
    .C(net414),
    .D(net882),
    .X(_00776_));
 sky130_fd_sc_hd__nor2_4 _09982_ (.A(_00774_),
    .B(_00776_),
    .Y(_00777_));
 sky130_fd_sc_hd__or3_4 _09983_ (.A(_00635_),
    .B(_00772_),
    .C(_00777_),
    .X(_00778_));
 sky130_fd_sc_hd__a22oi_4 _09984_ (.A1(net439),
    .A2(net843),
    .B1(net854),
    .B2(net430),
    .Y(_00779_));
 sky130_fd_sc_hd__and4_1 _09985_ (.A(net430),
    .B(net439),
    .C(net843),
    .D(net854),
    .X(_00780_));
 sky130_fd_sc_hd__nor2_2 _09986_ (.A(_00779_),
    .B(_00780_),
    .Y(_00781_));
 sky130_fd_sc_hd__nand2_4 _09987_ (.A(net449),
    .B(net833),
    .Y(_00782_));
 sky130_fd_sc_hd__xnor2_4 _09988_ (.A(_00781_),
    .B(_00782_),
    .Y(_00783_));
 sky130_fd_sc_hd__xnor2_4 _09989_ (.A(_00773_),
    .B(_00777_),
    .Y(_00784_));
 sky130_fd_sc_hd__nand2_2 _09990_ (.A(_00783_),
    .B(_00784_),
    .Y(_00785_));
 sky130_fd_sc_hd__a21oi_2 _09991_ (.A1(_00778_),
    .A2(_00785_),
    .B1(_00771_),
    .Y(_00786_));
 sky130_fd_sc_hd__a21o_1 _09992_ (.A1(_00778_),
    .A2(_00785_),
    .B1(_00771_),
    .X(_00787_));
 sky130_fd_sc_hd__o21ba_4 _09993_ (.A1(_00779_),
    .A2(_00782_),
    .B1_N(_00780_),
    .X(_00788_));
 sky130_fd_sc_hd__xnor2_4 _09994_ (.A(_00652_),
    .B(_00653_),
    .Y(_00789_));
 sky130_fd_sc_hd__nand2b_1 _09995_ (.A_N(_00788_),
    .B(_00789_),
    .Y(_00790_));
 sky130_fd_sc_hd__xnor2_4 _09996_ (.A(_00788_),
    .B(_00789_),
    .Y(_00791_));
 sky130_fd_sc_hd__and4_1 _09997_ (.A(net457),
    .B(net467),
    .C(net815),
    .D(net826),
    .X(_00792_));
 sky130_fd_sc_hd__nand2_4 _09998_ (.A(net475),
    .B(net806),
    .Y(_00793_));
 sky130_fd_sc_hd__a22oi_4 _09999_ (.A1(net467),
    .A2(net815),
    .B1(net826),
    .B2(net457),
    .Y(_00794_));
 sky130_fd_sc_hd__nor2_2 _10000_ (.A(_00792_),
    .B(_00794_),
    .Y(_00795_));
 sky130_fd_sc_hd__o21ba_4 _10001_ (.A1(_00793_),
    .A2(_00794_),
    .B1_N(_00792_),
    .X(_00796_));
 sky130_fd_sc_hd__nand2b_1 _10002_ (.A_N(_00796_),
    .B(_00791_),
    .Y(_00797_));
 sky130_fd_sc_hd__xnor2_4 _10003_ (.A(_00791_),
    .B(_00796_),
    .Y(_00798_));
 sky130_fd_sc_hd__nand3_2 _10004_ (.A(_00771_),
    .B(_00778_),
    .C(_00785_),
    .Y(_00799_));
 sky130_fd_sc_hd__and3_4 _10005_ (.A(_00787_),
    .B(_00798_),
    .C(_00799_),
    .X(_00800_));
 sky130_fd_sc_hd__o211a_1 _10006_ (.A1(_00786_),
    .A2(_00800_),
    .B1(_00659_),
    .C1(_00770_),
    .X(_00801_));
 sky130_fd_sc_hd__xnor2_2 _10007_ (.A(_00673_),
    .B(_00675_),
    .Y(_00802_));
 sky130_fd_sc_hd__a21o_1 _10008_ (.A1(_00790_),
    .A2(_00797_),
    .B1(_00802_),
    .X(_00803_));
 sky130_fd_sc_hd__nand3_1 _10009_ (.A(_00790_),
    .B(_00797_),
    .C(_00802_),
    .Y(_00804_));
 sky130_fd_sc_hd__nand2_1 _10010_ (.A(_00803_),
    .B(_00804_),
    .Y(_00805_));
 sky130_fd_sc_hd__o2bb2a_1 _10011_ (.A1_N(net502),
    .A2_N(net759),
    .B1(_00668_),
    .B2(_00669_),
    .X(_00806_));
 sky130_fd_sc_hd__nor2_2 _10012_ (.A(_00670_),
    .B(_00806_),
    .Y(_00807_));
 sky130_fd_sc_hd__nand2_4 _10013_ (.A(net499),
    .B(net793),
    .Y(_00808_));
 sky130_fd_sc_hd__and4_2 _10014_ (.A(net489),
    .B(net499),
    .C(net780),
    .D(net794),
    .X(_00809_));
 sky130_fd_sc_hd__a22oi_2 _10015_ (.A1(net499),
    .A2(net780),
    .B1(net794),
    .B2(net489),
    .Y(_00810_));
 sky130_fd_sc_hd__and4bb_2 _10016_ (.A_N(_00809_),
    .B_N(_00810_),
    .C(net506),
    .D(net770),
    .X(_00811_));
 sky130_fd_sc_hd__nor2_4 _10017_ (.A(_00809_),
    .B(_00811_),
    .Y(_00812_));
 sky130_fd_sc_hd__or3_1 _10018_ (.A(_00670_),
    .B(_00806_),
    .C(_00812_),
    .X(_00813_));
 sky130_fd_sc_hd__xnor2_4 _10019_ (.A(_00807_),
    .B(_00812_),
    .Y(_00814_));
 sky130_fd_sc_hd__o2bb2a_1 _10020_ (.A1_N(net531),
    .A2_N(net731),
    .B1(_00687_),
    .B2(_00688_),
    .X(_00815_));
 sky130_fd_sc_hd__nor2_2 _10021_ (.A(_00689_),
    .B(_00815_),
    .Y(_00816_));
 sky130_fd_sc_hd__nand2_1 _10022_ (.A(_00814_),
    .B(_00816_),
    .Y(_00817_));
 sky130_fd_sc_hd__nand3_1 _10023_ (.A(_00805_),
    .B(_00813_),
    .C(_00817_),
    .Y(_00818_));
 sky130_fd_sc_hd__a21o_2 _10024_ (.A1(_00813_),
    .A2(_00817_),
    .B1(_00805_),
    .X(_00819_));
 sky130_fd_sc_hd__a211oi_1 _10025_ (.A1(_00659_),
    .A2(_00770_),
    .B1(_00786_),
    .C1(_00800_),
    .Y(_00820_));
 sky130_fd_sc_hd__a211o_1 _10026_ (.A1(_00659_),
    .A2(_00770_),
    .B1(_00786_),
    .C1(_00800_),
    .X(_00821_));
 sky130_fd_sc_hd__and4b_4 _10027_ (.A_N(_00801_),
    .B(_00818_),
    .C(_00819_),
    .D(_00821_),
    .X(_00822_));
 sky130_fd_sc_hd__nor2_2 _10028_ (.A(_00801_),
    .B(_00822_),
    .Y(_00823_));
 sky130_fd_sc_hd__or3_1 _10029_ (.A(_00680_),
    .B(_00769_),
    .C(_00823_),
    .X(_00824_));
 sky130_fd_sc_hd__a21oi_2 _10030_ (.A1(_00699_),
    .A2(_00701_),
    .B1(_00703_),
    .Y(_00825_));
 sky130_fd_sc_hd__a211oi_2 _10031_ (.A1(_00803_),
    .A2(_00819_),
    .B1(_00825_),
    .C1(_00704_),
    .Y(_00826_));
 sky130_fd_sc_hd__o211a_1 _10032_ (.A1(_00704_),
    .A2(_00825_),
    .B1(_00819_),
    .C1(_00803_),
    .X(_00827_));
 sky130_fd_sc_hd__nor2_2 _10033_ (.A(_00826_),
    .B(_00827_),
    .Y(_00828_));
 sky130_fd_sc_hd__or3_1 _10034_ (.A(_00694_),
    .B(_00696_),
    .C(_00697_),
    .X(_00829_));
 sky130_fd_sc_hd__nand2_1 _10035_ (.A(_00698_),
    .B(_00829_),
    .Y(_00830_));
 sky130_fd_sc_hd__and4_2 _10036_ (.A(net514),
    .B(net521),
    .C(net748),
    .D(net759),
    .X(_00831_));
 sky130_fd_sc_hd__a22oi_2 _10037_ (.A1(net521),
    .A2(net748),
    .B1(net759),
    .B2(net514),
    .Y(_00832_));
 sky130_fd_sc_hd__and4bb_2 _10038_ (.A_N(_00831_),
    .B_N(_00832_),
    .C(net531),
    .D(net740),
    .X(_00833_));
 sky130_fd_sc_hd__nor2_4 _10039_ (.A(_00831_),
    .B(_00833_),
    .Y(_00834_));
 sky130_fd_sc_hd__o2bb2a_1 _10040_ (.A1_N(net574),
    .A2_N(net705),
    .B1(_00694_),
    .B2(_00695_),
    .X(_00835_));
 sky130_fd_sc_hd__nor2_2 _10041_ (.A(_00696_),
    .B(_00835_),
    .Y(_00836_));
 sky130_fd_sc_hd__or3_2 _10042_ (.A(_00696_),
    .B(_00834_),
    .C(_00835_),
    .X(_00837_));
 sky130_fd_sc_hd__and4_2 _10043_ (.A(net543),
    .B(net557),
    .C(net722),
    .D(net731),
    .X(_00838_));
 sky130_fd_sc_hd__a22oi_2 _10044_ (.A1(net557),
    .A2(net722),
    .B1(net731),
    .B2(net543),
    .Y(_00839_));
 sky130_fd_sc_hd__and4bb_4 _10045_ (.A_N(_00838_),
    .B_N(_00839_),
    .C(net574),
    .D(net713),
    .X(_00840_));
 sky130_fd_sc_hd__xnor2_4 _10046_ (.A(_00834_),
    .B(_00836_),
    .Y(_00841_));
 sky130_fd_sc_hd__o21ai_4 _10047_ (.A1(_00838_),
    .A2(_00840_),
    .B1(_00841_),
    .Y(_00842_));
 sky130_fd_sc_hd__a21o_2 _10048_ (.A1(_00837_),
    .A2(_00842_),
    .B1(_00830_),
    .X(_00843_));
 sky130_fd_sc_hd__inv_2 _10049_ (.A(_00843_),
    .Y(_00844_));
 sky130_fd_sc_hd__nand3_2 _10050_ (.A(_00830_),
    .B(_00837_),
    .C(_00842_),
    .Y(_00845_));
 sky130_fd_sc_hd__o21ai_1 _10051_ (.A1(_00577_),
    .A2(_00719_),
    .B1(_00724_),
    .Y(_00846_));
 sky130_fd_sc_hd__and2_2 _10052_ (.A(_00725_),
    .B(_00846_),
    .X(_00847_));
 sky130_fd_sc_hd__and3_4 _10053_ (.A(_00843_),
    .B(_00845_),
    .C(_00847_),
    .X(_00848_));
 sky130_fd_sc_hd__nor2_4 _10054_ (.A(_00844_),
    .B(_00848_),
    .Y(_00849_));
 sky130_fd_sc_hd__xnor2_4 _10055_ (.A(_00828_),
    .B(_00849_),
    .Y(_00850_));
 sky130_fd_sc_hd__o21ai_4 _10056_ (.A1(_00680_),
    .A2(_00769_),
    .B1(_00823_),
    .Y(_00851_));
 sky130_fd_sc_hd__and3_1 _10057_ (.A(_00824_),
    .B(_00850_),
    .C(_00851_),
    .X(_00852_));
 sky130_fd_sc_hd__a21boi_4 _10058_ (.A1(_00850_),
    .A2(_00851_),
    .B1_N(_00824_),
    .Y(_00853_));
 sky130_fd_sc_hd__nor3_4 _10059_ (.A(_00711_),
    .B(_00768_),
    .C(_00853_),
    .Y(_00854_));
 sky130_fd_sc_hd__inv_2 _10060_ (.A(_00854_),
    .Y(_00855_));
 sky130_fd_sc_hd__xnor2_2 _10061_ (.A(_00742_),
    .B(_00743_),
    .Y(_00856_));
 sky130_fd_sc_hd__and3_2 _10062_ (.A(net381),
    .B(net911),
    .C(_00591_),
    .X(_00857_));
 sky130_fd_sc_hd__o2bb2a_1 _10063_ (.A1_N(net382),
    .A2_N(net893),
    .B1(_00737_),
    .B2(_00738_),
    .X(_00858_));
 sky130_fd_sc_hd__nor2_1 _10064_ (.A(_00739_),
    .B(_00858_),
    .Y(_00859_));
 sky130_fd_sc_hd__and2_2 _10065_ (.A(_00857_),
    .B(_00859_),
    .X(_00860_));
 sky130_fd_sc_hd__xor2_1 _10066_ (.A(_00857_),
    .B(_00859_),
    .X(_00861_));
 sky130_fd_sc_hd__and3_2 _10067_ (.A(net390),
    .B(net882),
    .C(_00861_),
    .X(_00862_));
 sky130_fd_sc_hd__o21ai_4 _10068_ (.A1(_00860_),
    .A2(_00862_),
    .B1(_00856_),
    .Y(_00863_));
 sky130_fd_sc_hd__or3_1 _10069_ (.A(_00856_),
    .B(_00860_),
    .C(_00862_),
    .X(_00864_));
 sky130_fd_sc_hd__and2_2 _10070_ (.A(_00863_),
    .B(_00864_),
    .X(_00865_));
 sky130_fd_sc_hd__nand2_1 _10071_ (.A(net398),
    .B(net863),
    .Y(_00866_));
 sky130_fd_sc_hd__nand3_2 _10072_ (.A(net398),
    .B(net863),
    .C(_00865_),
    .Y(_00867_));
 sky130_fd_sc_hd__xor2_2 _10073_ (.A(_00865_),
    .B(_00866_),
    .X(_00868_));
 sky130_fd_sc_hd__nand2_1 _10074_ (.A(_00296_),
    .B(_00725_),
    .Y(_00869_));
 sky130_fd_sc_hd__nand2_1 _10075_ (.A(_00726_),
    .B(_00869_),
    .Y(_00870_));
 sky130_fd_sc_hd__nor2_2 _10076_ (.A(_00868_),
    .B(_00870_),
    .Y(_00871_));
 sky130_fd_sc_hd__o21bai_2 _10077_ (.A1(_00827_),
    .A2(_00849_),
    .B1_N(_00826_),
    .Y(_00872_));
 sky130_fd_sc_hd__xor2_2 _10078_ (.A(_00731_),
    .B(_00748_),
    .X(_00873_));
 sky130_fd_sc_hd__nand2_2 _10079_ (.A(_00872_),
    .B(_00873_),
    .Y(_00874_));
 sky130_fd_sc_hd__or2_1 _10080_ (.A(_00872_),
    .B(_00873_),
    .X(_00875_));
 sky130_fd_sc_hd__and2_1 _10081_ (.A(_00874_),
    .B(_00875_),
    .X(_00876_));
 sky130_fd_sc_hd__nand2_2 _10082_ (.A(_00871_),
    .B(_00876_),
    .Y(_00877_));
 sky130_fd_sc_hd__or2_1 _10083_ (.A(_00871_),
    .B(_00876_),
    .X(_00878_));
 sky130_fd_sc_hd__nand2_2 _10084_ (.A(_00877_),
    .B(_00878_),
    .Y(_00879_));
 sky130_fd_sc_hd__o21a_2 _10085_ (.A1(_00711_),
    .A2(_00768_),
    .B1(_00853_),
    .X(_00880_));
 sky130_fd_sc_hd__or3_4 _10086_ (.A(_00854_),
    .B(_00879_),
    .C(_00880_),
    .X(_00881_));
 sky130_fd_sc_hd__a211oi_4 _10087_ (.A1(_00855_),
    .A2(_00881_),
    .B1(_00754_),
    .C1(_00767_),
    .Y(_00882_));
 sky130_fd_sc_hd__o211a_2 _10088_ (.A1(_00754_),
    .A2(_00767_),
    .B1(_00855_),
    .C1(_00881_),
    .X(_00883_));
 sky130_fd_sc_hd__a211oi_4 _10089_ (.A1(_00874_),
    .A2(_00877_),
    .B1(_00882_),
    .C1(_00883_),
    .Y(_00884_));
 sky130_fd_sc_hd__nor2_2 _10090_ (.A(_00882_),
    .B(_00884_),
    .Y(_00885_));
 sky130_fd_sc_hd__nor3_4 _10091_ (.A(_00758_),
    .B(_00766_),
    .C(_00885_),
    .Y(_00886_));
 sky130_fd_sc_hd__o21a_2 _10092_ (.A1(_00758_),
    .A2(_00766_),
    .B1(_00885_),
    .X(_00887_));
 sky130_fd_sc_hd__a211oi_4 _10093_ (.A1(_00599_),
    .A2(_00602_),
    .B1(_00886_),
    .C1(_00887_),
    .Y(_00888_));
 sky130_fd_sc_hd__nor2_2 _10094_ (.A(_00886_),
    .B(_00888_),
    .Y(_00889_));
 sky130_fd_sc_hd__or2_1 _10095_ (.A(_00765_),
    .B(_00889_),
    .X(_00890_));
 sky130_fd_sc_hd__o21ai_4 _10096_ (.A1(_00760_),
    .A2(_00762_),
    .B1(_00622_),
    .Y(_00891_));
 sky130_fd_sc_hd__nand2_1 _10097_ (.A(_00765_),
    .B(_00889_),
    .Y(_00892_));
 sky130_fd_sc_hd__and2_4 _10098_ (.A(_00890_),
    .B(_00892_),
    .X(_00893_));
 sky130_fd_sc_hd__o211a_2 _10099_ (.A1(_00886_),
    .A2(_00887_),
    .B1(_00599_),
    .C1(_00602_),
    .X(_00894_));
 sky130_fd_sc_hd__o211a_1 _10100_ (.A1(_00882_),
    .A2(_00883_),
    .B1(_00874_),
    .C1(_00877_),
    .X(_00895_));
 sky130_fd_sc_hd__nor2_4 _10101_ (.A(_00884_),
    .B(_00895_),
    .Y(_00896_));
 sky130_fd_sc_hd__o21ai_4 _10102_ (.A1(_00854_),
    .A2(_00880_),
    .B1(_00879_),
    .Y(_00897_));
 sky130_fd_sc_hd__a21oi_1 _10103_ (.A1(_00824_),
    .A2(_00851_),
    .B1(_00850_),
    .Y(_00898_));
 sky130_fd_sc_hd__o2bb2a_2 _10104_ (.A1_N(_00818_),
    .A2_N(_00819_),
    .B1(_00820_),
    .B2(_00801_),
    .X(_00899_));
 sky130_fd_sc_hd__a21oi_4 _10105_ (.A1(_00787_),
    .A2(_00799_),
    .B1(_00798_),
    .Y(_00900_));
 sky130_fd_sc_hd__xnor2_4 _10106_ (.A(_00783_),
    .B(_00784_),
    .Y(_00901_));
 sky130_fd_sc_hd__o2bb2a_1 _10107_ (.A1_N(net414),
    .A2_N(net882),
    .B1(_00774_),
    .B2(_00775_),
    .X(_00902_));
 sky130_fd_sc_hd__nor2_2 _10108_ (.A(_00776_),
    .B(_00902_),
    .Y(_00903_));
 sky130_fd_sc_hd__and4_2 _10109_ (.A(net406),
    .B(net422),
    .C(net882),
    .D(net904),
    .X(_00904_));
 sky130_fd_sc_hd__a22oi_2 _10110_ (.A1(net422),
    .A2(net882),
    .B1(net904),
    .B2(net406),
    .Y(_00905_));
 sky130_fd_sc_hd__and4bb_4 _10111_ (.A_N(_00904_),
    .B_N(_00905_),
    .C(net414),
    .D(net894),
    .X(_00906_));
 sky130_fd_sc_hd__nor2_4 _10112_ (.A(_00904_),
    .B(_00906_),
    .Y(_00907_));
 sky130_fd_sc_hd__or3_4 _10113_ (.A(_00776_),
    .B(_00902_),
    .C(_00907_),
    .X(_00908_));
 sky130_fd_sc_hd__a22oi_4 _10114_ (.A1(net439),
    .A2(net854),
    .B1(net863),
    .B2(net430),
    .Y(_00909_));
 sky130_fd_sc_hd__and4_1 _10115_ (.A(net430),
    .B(net439),
    .C(net854),
    .D(net863),
    .X(_00910_));
 sky130_fd_sc_hd__nor2_2 _10116_ (.A(_00909_),
    .B(_00910_),
    .Y(_00911_));
 sky130_fd_sc_hd__nand2_4 _10117_ (.A(net447),
    .B(net843),
    .Y(_00912_));
 sky130_fd_sc_hd__xnor2_4 _10118_ (.A(_00911_),
    .B(_00912_),
    .Y(_00913_));
 sky130_fd_sc_hd__xnor2_4 _10119_ (.A(_00903_),
    .B(_00907_),
    .Y(_00914_));
 sky130_fd_sc_hd__nand2_2 _10120_ (.A(_00913_),
    .B(_00914_),
    .Y(_00915_));
 sky130_fd_sc_hd__a21o_4 _10121_ (.A1(_00908_),
    .A2(_00915_),
    .B1(_00901_),
    .X(_00916_));
 sky130_fd_sc_hd__o21ba_4 _10122_ (.A1(_00909_),
    .A2(_00912_),
    .B1_N(_00910_),
    .X(_00917_));
 sky130_fd_sc_hd__xnor2_4 _10123_ (.A(_00793_),
    .B(_00795_),
    .Y(_00918_));
 sky130_fd_sc_hd__nand2b_2 _10124_ (.A_N(_00917_),
    .B(_00918_),
    .Y(_00919_));
 sky130_fd_sc_hd__xnor2_4 _10125_ (.A(_00917_),
    .B(_00918_),
    .Y(_00920_));
 sky130_fd_sc_hd__and4_1 _10126_ (.A(net457),
    .B(net467),
    .C(net826),
    .D(net833),
    .X(_00921_));
 sky130_fd_sc_hd__a22oi_4 _10127_ (.A1(net467),
    .A2(net826),
    .B1(net833),
    .B2(net457),
    .Y(_00922_));
 sky130_fd_sc_hd__nor2_2 _10128_ (.A(_00921_),
    .B(_00922_),
    .Y(_00923_));
 sky130_fd_sc_hd__nand2_4 _10129_ (.A(net475),
    .B(net815),
    .Y(_00924_));
 sky130_fd_sc_hd__o21ba_1 _10130_ (.A1(_00922_),
    .A2(_00924_),
    .B1_N(_00921_),
    .X(_00925_));
 sky130_fd_sc_hd__nand2b_2 _10131_ (.A_N(_00925_),
    .B(_00920_),
    .Y(_00926_));
 sky130_fd_sc_hd__xnor2_2 _10132_ (.A(_00920_),
    .B(_00925_),
    .Y(_00927_));
 sky130_fd_sc_hd__nand3_4 _10133_ (.A(_00901_),
    .B(_00908_),
    .C(_00915_),
    .Y(_00928_));
 sky130_fd_sc_hd__nand3_4 _10134_ (.A(_00916_),
    .B(_00927_),
    .C(_00928_),
    .Y(_00929_));
 sky130_fd_sc_hd__a211o_4 _10135_ (.A1(_00916_),
    .A2(_00929_),
    .B1(_00800_),
    .C1(_00900_),
    .X(_00930_));
 sky130_fd_sc_hd__xnor2_2 _10136_ (.A(_00814_),
    .B(_00816_),
    .Y(_00931_));
 sky130_fd_sc_hd__a21o_4 _10137_ (.A1(_00919_),
    .A2(_00926_),
    .B1(_00931_),
    .X(_00932_));
 sky130_fd_sc_hd__nand3_2 _10138_ (.A(_00919_),
    .B(_00926_),
    .C(_00931_),
    .Y(_00933_));
 sky130_fd_sc_hd__o2bb2a_1 _10139_ (.A1_N(net506),
    .A2_N(net770),
    .B1(_00809_),
    .B2(_00810_),
    .X(_00934_));
 sky130_fd_sc_hd__nor2_2 _10140_ (.A(_00811_),
    .B(_00934_),
    .Y(_00935_));
 sky130_fd_sc_hd__and2_4 _10141_ (.A(net489),
    .B(net806),
    .X(_00936_));
 sky130_fd_sc_hd__nand2_4 _10142_ (.A(net489),
    .B(net806),
    .Y(_00937_));
 sky130_fd_sc_hd__nor2_2 _10143_ (.A(_00808_),
    .B(_00937_),
    .Y(_00938_));
 sky130_fd_sc_hd__nand2_1 _10144_ (.A(net506),
    .B(net780),
    .Y(_00939_));
 sky130_fd_sc_hd__xnor2_4 _10145_ (.A(_00808_),
    .B(_00936_),
    .Y(_00940_));
 sky130_fd_sc_hd__and3_1 _10146_ (.A(net506),
    .B(net780),
    .C(_00940_),
    .X(_00941_));
 sky130_fd_sc_hd__o21a_4 _10147_ (.A1(_00938_),
    .A2(_00941_),
    .B1(_00935_),
    .X(_00942_));
 sky130_fd_sc_hd__nor3_2 _10148_ (.A(_00935_),
    .B(_00938_),
    .C(_00941_),
    .Y(_00943_));
 sky130_fd_sc_hd__nor2_4 _10149_ (.A(_00942_),
    .B(_00943_),
    .Y(_00944_));
 sky130_fd_sc_hd__o2bb2a_1 _10150_ (.A1_N(net531),
    .A2_N(net740),
    .B1(_00831_),
    .B2(_00832_),
    .X(_00945_));
 sky130_fd_sc_hd__nor2_2 _10151_ (.A(_00833_),
    .B(_00945_),
    .Y(_00946_));
 sky130_fd_sc_hd__and2_2 _10152_ (.A(_00944_),
    .B(_00946_),
    .X(_00947_));
 sky130_fd_sc_hd__o211ai_4 _10153_ (.A1(_00942_),
    .A2(_00947_),
    .B1(_00932_),
    .C1(_00933_),
    .Y(_00948_));
 sky130_fd_sc_hd__a211o_1 _10154_ (.A1(_00932_),
    .A2(_00933_),
    .B1(_00942_),
    .C1(_00947_),
    .X(_00949_));
 sky130_fd_sc_hd__nand2_1 _10155_ (.A(_00948_),
    .B(_00949_),
    .Y(_00950_));
 sky130_fd_sc_hd__o211ai_4 _10156_ (.A1(_00800_),
    .A2(_00900_),
    .B1(_00916_),
    .C1(_00929_),
    .Y(_00951_));
 sky130_fd_sc_hd__nand3b_4 _10157_ (.A_N(_00950_),
    .B(_00951_),
    .C(_00930_),
    .Y(_00952_));
 sky130_fd_sc_hd__a211oi_4 _10158_ (.A1(_00930_),
    .A2(_00952_),
    .B1(_00822_),
    .C1(_00899_),
    .Y(_00953_));
 sky130_fd_sc_hd__a21oi_4 _10159_ (.A1(_00843_),
    .A2(_00845_),
    .B1(_00847_),
    .Y(_00954_));
 sky130_fd_sc_hd__a211oi_4 _10160_ (.A1(_00932_),
    .A2(_00948_),
    .B1(_00954_),
    .C1(_00848_),
    .Y(_00955_));
 sky130_fd_sc_hd__o211a_2 _10161_ (.A1(_00848_),
    .A2(_00954_),
    .B1(_00948_),
    .C1(_00932_),
    .X(_00956_));
 sky130_fd_sc_hd__or3_1 _10162_ (.A(_00838_),
    .B(_00840_),
    .C(_00841_),
    .X(_00957_));
 sky130_fd_sc_hd__nand2_2 _10163_ (.A(_00842_),
    .B(_00957_),
    .Y(_00958_));
 sky130_fd_sc_hd__and4_1 _10164_ (.A(net514),
    .B(net521),
    .C(net757),
    .D(net768),
    .X(_00959_));
 sky130_fd_sc_hd__a22oi_2 _10165_ (.A1(net521),
    .A2(net757),
    .B1(net768),
    .B2(net514),
    .Y(_00960_));
 sky130_fd_sc_hd__and4bb_1 _10166_ (.A_N(_00959_),
    .B_N(_00960_),
    .C(net531),
    .D(net748),
    .X(_00961_));
 sky130_fd_sc_hd__nor2_2 _10167_ (.A(_00959_),
    .B(_00961_),
    .Y(_00962_));
 sky130_fd_sc_hd__o2bb2a_1 _10168_ (.A1_N(net574),
    .A2_N(net713),
    .B1(_00838_),
    .B2(_00839_),
    .X(_00963_));
 sky130_fd_sc_hd__nor2_1 _10169_ (.A(_00840_),
    .B(_00963_),
    .Y(_00964_));
 sky130_fd_sc_hd__or3_4 _10170_ (.A(_00840_),
    .B(_00962_),
    .C(_00963_),
    .X(_00965_));
 sky130_fd_sc_hd__and4_2 _10171_ (.A(net543),
    .B(net557),
    .C(net731),
    .D(net740),
    .X(_00966_));
 sky130_fd_sc_hd__a22oi_2 _10172_ (.A1(net557),
    .A2(net731),
    .B1(net740),
    .B2(net543),
    .Y(_00967_));
 sky130_fd_sc_hd__and4bb_4 _10173_ (.A_N(_00966_),
    .B_N(_00967_),
    .C(net574),
    .D(net722),
    .X(_00968_));
 sky130_fd_sc_hd__xnor2_2 _10174_ (.A(_00962_),
    .B(_00964_),
    .Y(_00969_));
 sky130_fd_sc_hd__o21ai_4 _10175_ (.A1(_00966_),
    .A2(_00968_),
    .B1(_00969_),
    .Y(_00970_));
 sky130_fd_sc_hd__a21o_4 _10176_ (.A1(_00965_),
    .A2(_00970_),
    .B1(_00958_),
    .X(_00971_));
 sky130_fd_sc_hd__nand3_4 _10177_ (.A(_00958_),
    .B(_00965_),
    .C(_00970_),
    .Y(_00972_));
 sky130_fd_sc_hd__o2bb2a_1 _10178_ (.A1_N(\ApproximateM_inst.lob_16.lob2.genblk1[1].genblk1.mux.sel ),
    .A2_N(net687),
    .B1(_00721_),
    .B2(_00722_),
    .X(_00973_));
 sky130_fd_sc_hd__and2_2 _10179_ (.A(net609),
    .B(net704),
    .X(_00974_));
 sky130_fd_sc_hd__and3_1 _10180_ (.A(net582),
    .B(net688),
    .C(_00974_),
    .X(_00975_));
 sky130_fd_sc_hd__a21oi_1 _10181_ (.A1(net582),
    .A2(net704),
    .B1(_00574_),
    .Y(_00976_));
 sky130_fd_sc_hd__and4bb_2 _10182_ (.A_N(_00975_),
    .B_N(_00976_),
    .C(net594),
    .D(net696),
    .X(_00977_));
 sky130_fd_sc_hd__nor2_1 _10183_ (.A(_00975_),
    .B(_00977_),
    .Y(_00978_));
 sky130_fd_sc_hd__or3_4 _10184_ (.A(_00723_),
    .B(_00973_),
    .C(_00978_),
    .X(_00979_));
 sky130_fd_sc_hd__o21ai_1 _10185_ (.A1(_00723_),
    .A2(_00973_),
    .B1(_00978_),
    .Y(_00980_));
 sky130_fd_sc_hd__and2_4 _10186_ (.A(_00979_),
    .B(_00980_),
    .X(_00981_));
 sky130_fd_sc_hd__and3_2 _10187_ (.A(_00971_),
    .B(_00972_),
    .C(_00981_),
    .X(_00982_));
 sky130_fd_sc_hd__nand3_2 _10188_ (.A(_00971_),
    .B(_00972_),
    .C(_00981_),
    .Y(_00983_));
 sky130_fd_sc_hd__o211a_2 _10189_ (.A1(_00955_),
    .A2(_00956_),
    .B1(_00971_),
    .C1(_00983_),
    .X(_00984_));
 sky130_fd_sc_hd__a211oi_4 _10190_ (.A1(_00971_),
    .A2(_00983_),
    .B1(_00955_),
    .C1(_00956_),
    .Y(_00985_));
 sky130_fd_sc_hd__o211a_2 _10191_ (.A1(_00822_),
    .A2(_00899_),
    .B1(_00930_),
    .C1(_00952_),
    .X(_00986_));
 sky130_fd_sc_hd__nor4_4 _10192_ (.A(_00953_),
    .B(_00984_),
    .C(_00985_),
    .D(_00986_),
    .Y(_00987_));
 sky130_fd_sc_hd__nor2_1 _10193_ (.A(_00953_),
    .B(_00987_),
    .Y(_00988_));
 sky130_fd_sc_hd__nor3_1 _10194_ (.A(_00852_),
    .B(_00898_),
    .C(_00988_),
    .Y(_00989_));
 sky130_fd_sc_hd__nand2_4 _10195_ (.A(net390),
    .B(net893),
    .Y(_00990_));
 sky130_fd_sc_hd__a22oi_4 _10196_ (.A1(net381),
    .A2(net902),
    .B1(net911),
    .B2(net374),
    .Y(_00991_));
 sky130_fd_sc_hd__nor2_2 _10197_ (.A(_00857_),
    .B(_00991_),
    .Y(_00992_));
 sky130_fd_sc_hd__or3_2 _10198_ (.A(_00857_),
    .B(_00990_),
    .C(_00991_),
    .X(_00993_));
 sky130_fd_sc_hd__a21oi_1 _10199_ (.A1(net390),
    .A2(net882),
    .B1(_00861_),
    .Y(_00994_));
 sky130_fd_sc_hd__nor2_2 _10200_ (.A(_00862_),
    .B(_00994_),
    .Y(_00995_));
 sky130_fd_sc_hd__and2b_1 _10201_ (.A_N(_00993_),
    .B(_00995_),
    .X(_00996_));
 sky130_fd_sc_hd__xnor2_2 _10202_ (.A(_00993_),
    .B(_00995_),
    .Y(_00997_));
 sky130_fd_sc_hd__and3_2 _10203_ (.A(net397),
    .B(net872),
    .C(_00997_),
    .X(_00998_));
 sky130_fd_sc_hd__a21oi_2 _10204_ (.A1(net397),
    .A2(net872),
    .B1(_00997_),
    .Y(_00999_));
 sky130_fd_sc_hd__nor2_4 _10205_ (.A(_00998_),
    .B(_00999_),
    .Y(_01000_));
 sky130_fd_sc_hd__and2b_1 _10206_ (.A_N(_00979_),
    .B(_01000_),
    .X(_01001_));
 sky130_fd_sc_hd__nor2_2 _10207_ (.A(_00955_),
    .B(_00985_),
    .Y(_01002_));
 sky130_fd_sc_hd__and2_1 _10208_ (.A(_00868_),
    .B(_00870_),
    .X(_01003_));
 sky130_fd_sc_hd__nor2_1 _10209_ (.A(_00871_),
    .B(_01003_),
    .Y(_01004_));
 sky130_fd_sc_hd__xnor2_2 _10210_ (.A(_01002_),
    .B(_01004_),
    .Y(_01005_));
 sky130_fd_sc_hd__nand2_1 _10211_ (.A(_01001_),
    .B(_01005_),
    .Y(_01006_));
 sky130_fd_sc_hd__xnor2_1 _10212_ (.A(_01001_),
    .B(_01005_),
    .Y(_01007_));
 sky130_fd_sc_hd__o21a_1 _10213_ (.A1(_00852_),
    .A2(_00898_),
    .B1(_00988_),
    .X(_01008_));
 sky130_fd_sc_hd__or3_2 _10214_ (.A(_00989_),
    .B(_01007_),
    .C(_01008_),
    .X(_01009_));
 sky130_fd_sc_hd__nand2b_2 _10215_ (.A_N(_00989_),
    .B(_01009_),
    .Y(_01010_));
 sky130_fd_sc_hd__and3_2 _10216_ (.A(_00881_),
    .B(_00897_),
    .C(_01010_),
    .X(_01011_));
 sky130_fd_sc_hd__o31a_2 _10217_ (.A1(_00871_),
    .A2(_01002_),
    .A3(_01003_),
    .B1(_01006_),
    .X(_01012_));
 sky130_fd_sc_hd__a21oi_4 _10218_ (.A1(_00881_),
    .A2(_00897_),
    .B1(_01010_),
    .Y(_01013_));
 sky130_fd_sc_hd__or3_4 _10219_ (.A(_01011_),
    .B(_01012_),
    .C(_01013_),
    .X(_01014_));
 sky130_fd_sc_hd__and2b_2 _10220_ (.A_N(_01011_),
    .B(_01014_),
    .X(_01015_));
 sky130_fd_sc_hd__and2b_1 _10221_ (.A_N(_01015_),
    .B(_00896_),
    .X(_01016_));
 sky130_fd_sc_hd__a31o_4 _10222_ (.A1(net398),
    .A2(net854),
    .A3(_00747_),
    .B1(_00745_),
    .X(_01017_));
 sky130_fd_sc_hd__xnor2_4 _10223_ (.A(_00896_),
    .B(_01015_),
    .Y(_01018_));
 sky130_fd_sc_hd__a21oi_2 _10224_ (.A1(_01017_),
    .A2(_01018_),
    .B1(_01016_),
    .Y(_01019_));
 sky130_fd_sc_hd__o21ai_4 _10225_ (.A1(_00888_),
    .A2(_00894_),
    .B1(_01019_),
    .Y(_01020_));
 sky130_fd_sc_hd__xnor2_4 _10226_ (.A(_01017_),
    .B(_01018_),
    .Y(_01021_));
 sky130_fd_sc_hd__o21ai_4 _10227_ (.A1(_01011_),
    .A2(_01013_),
    .B1(_01012_),
    .Y(_01022_));
 sky130_fd_sc_hd__o21ai_1 _10228_ (.A1(_00989_),
    .A2(_01008_),
    .B1(_01007_),
    .Y(_01023_));
 sky130_fd_sc_hd__o22a_2 _10229_ (.A1(_00984_),
    .A2(_00985_),
    .B1(_00986_),
    .B2(_00953_),
    .X(_01024_));
 sky130_fd_sc_hd__a21bo_2 _10230_ (.A1(_00930_),
    .A2(_00951_),
    .B1_N(_00950_),
    .X(_01025_));
 sky130_fd_sc_hd__a21o_1 _10231_ (.A1(_00916_),
    .A2(_00928_),
    .B1(_00927_),
    .X(_01026_));
 sky130_fd_sc_hd__xnor2_4 _10232_ (.A(_00913_),
    .B(_00914_),
    .Y(_01027_));
 sky130_fd_sc_hd__o2bb2a_1 _10233_ (.A1_N(net414),
    .A2_N(net894),
    .B1(_00904_),
    .B2(_00905_),
    .X(_01028_));
 sky130_fd_sc_hd__nor2_4 _10234_ (.A(_00906_),
    .B(_01028_),
    .Y(_01029_));
 sky130_fd_sc_hd__nand2_4 _10235_ (.A(net422),
    .B(net913),
    .Y(_01030_));
 sky130_fd_sc_hd__and4_1 _10236_ (.A(net406),
    .B(net422),
    .C(net894),
    .D(net913),
    .X(_01031_));
 sky130_fd_sc_hd__a22o_1 _10237_ (.A1(net422),
    .A2(net894),
    .B1(net913),
    .B2(net406),
    .X(_01032_));
 sky130_fd_sc_hd__nand2_1 _10238_ (.A(net414),
    .B(net904),
    .Y(_01033_));
 sky130_fd_sc_hd__a31o_4 _10239_ (.A1(net414),
    .A2(net904),
    .A3(_01032_),
    .B1(_01031_),
    .X(_01034_));
 sky130_fd_sc_hd__nand2_2 _10240_ (.A(_01029_),
    .B(_01034_),
    .Y(_01035_));
 sky130_fd_sc_hd__and4_1 _10241_ (.A(net430),
    .B(net439),
    .C(net863),
    .D(net872),
    .X(_01036_));
 sky130_fd_sc_hd__a22oi_4 _10242_ (.A1(net439),
    .A2(net863),
    .B1(net872),
    .B2(net430),
    .Y(_01037_));
 sky130_fd_sc_hd__nor2_2 _10243_ (.A(_01036_),
    .B(_01037_),
    .Y(_01038_));
 sky130_fd_sc_hd__nand2_4 _10244_ (.A(net447),
    .B(net854),
    .Y(_01039_));
 sky130_fd_sc_hd__xnor2_4 _10245_ (.A(_01038_),
    .B(_01039_),
    .Y(_01040_));
 sky130_fd_sc_hd__xor2_4 _10246_ (.A(_01029_),
    .B(_01034_),
    .X(_01041_));
 sky130_fd_sc_hd__nand2_2 _10247_ (.A(_01040_),
    .B(_01041_),
    .Y(_01042_));
 sky130_fd_sc_hd__a21o_2 _10248_ (.A1(_01035_),
    .A2(_01042_),
    .B1(_01027_),
    .X(_01043_));
 sky130_fd_sc_hd__inv_2 _10249_ (.A(_01043_),
    .Y(_01044_));
 sky130_fd_sc_hd__o21ba_4 _10250_ (.A1(_01037_),
    .A2(_01039_),
    .B1_N(_01036_),
    .X(_01045_));
 sky130_fd_sc_hd__xnor2_4 _10251_ (.A(_00923_),
    .B(_00924_),
    .Y(_01046_));
 sky130_fd_sc_hd__nand2b_2 _10252_ (.A_N(_01045_),
    .B(_01046_),
    .Y(_01047_));
 sky130_fd_sc_hd__xnor2_4 _10253_ (.A(_01045_),
    .B(_01046_),
    .Y(_01048_));
 sky130_fd_sc_hd__and4_1 _10254_ (.A(net457),
    .B(net467),
    .C(net833),
    .D(net843),
    .X(_01049_));
 sky130_fd_sc_hd__nand2_2 _10255_ (.A(net475),
    .B(net825),
    .Y(_01050_));
 sky130_fd_sc_hd__a22oi_2 _10256_ (.A1(net467),
    .A2(net833),
    .B1(net843),
    .B2(net457),
    .Y(_01051_));
 sky130_fd_sc_hd__nor2_1 _10257_ (.A(_01049_),
    .B(_01051_),
    .Y(_01052_));
 sky130_fd_sc_hd__o21ba_2 _10258_ (.A1(_01050_),
    .A2(_01051_),
    .B1_N(_01049_),
    .X(_01053_));
 sky130_fd_sc_hd__nand2b_2 _10259_ (.A_N(_01053_),
    .B(_01048_),
    .Y(_01054_));
 sky130_fd_sc_hd__xnor2_4 _10260_ (.A(_01048_),
    .B(_01053_),
    .Y(_01055_));
 sky130_fd_sc_hd__nand3_4 _10261_ (.A(_01027_),
    .B(_01035_),
    .C(_01042_),
    .Y(_01056_));
 sky130_fd_sc_hd__and3_4 _10262_ (.A(_01043_),
    .B(_01055_),
    .C(_01056_),
    .X(_01057_));
 sky130_fd_sc_hd__o211a_2 _10263_ (.A1(_01044_),
    .A2(_01057_),
    .B1(_00929_),
    .C1(_01026_),
    .X(_01058_));
 sky130_fd_sc_hd__o211ai_2 _10264_ (.A1(_01044_),
    .A2(_01057_),
    .B1(_00929_),
    .C1(_01026_),
    .Y(_01059_));
 sky130_fd_sc_hd__xnor2_4 _10265_ (.A(_00944_),
    .B(_00946_),
    .Y(_01060_));
 sky130_fd_sc_hd__a21o_4 _10266_ (.A1(_01047_),
    .A2(_01054_),
    .B1(_01060_),
    .X(_01061_));
 sky130_fd_sc_hd__nand3_2 _10267_ (.A(_01047_),
    .B(_01054_),
    .C(_01060_),
    .Y(_01062_));
 sky130_fd_sc_hd__xnor2_2 _10268_ (.A(_00939_),
    .B(_00940_),
    .Y(_01063_));
 sky130_fd_sc_hd__and2_2 _10269_ (.A(net499),
    .B(net816),
    .X(_01064_));
 sky130_fd_sc_hd__nand2_1 _10270_ (.A(net499),
    .B(net816),
    .Y(_01065_));
 sky130_fd_sc_hd__nand2_2 _10271_ (.A(net506),
    .B(net791),
    .Y(_01066_));
 sky130_fd_sc_hd__a22o_1 _10272_ (.A1(net499),
    .A2(net805),
    .B1(net814),
    .B2(net489),
    .X(_01067_));
 sky130_fd_sc_hd__o21a_4 _10273_ (.A1(_00937_),
    .A2(_01065_),
    .B1(_01067_),
    .X(_01068_));
 sky130_fd_sc_hd__a32o_4 _10274_ (.A1(net506),
    .A2(net792),
    .A3(_01067_),
    .B1(_01064_),
    .B2(_00936_),
    .X(_01069_));
 sky130_fd_sc_hd__and2_2 _10275_ (.A(_01063_),
    .B(_01069_),
    .X(_01070_));
 sky130_fd_sc_hd__xor2_2 _10276_ (.A(_01063_),
    .B(_01069_),
    .X(_01071_));
 sky130_fd_sc_hd__o2bb2a_1 _10277_ (.A1_N(net531),
    .A2_N(net748),
    .B1(_00959_),
    .B2(_00960_),
    .X(_01072_));
 sky130_fd_sc_hd__nor2_1 _10278_ (.A(_00961_),
    .B(_01072_),
    .Y(_01073_));
 sky130_fd_sc_hd__and2_2 _10279_ (.A(_01071_),
    .B(_01073_),
    .X(_01074_));
 sky130_fd_sc_hd__a211o_1 _10280_ (.A1(_01061_),
    .A2(_01062_),
    .B1(_01070_),
    .C1(_01074_),
    .X(_01075_));
 sky130_fd_sc_hd__o211ai_4 _10281_ (.A1(_01070_),
    .A2(_01074_),
    .B1(_01061_),
    .C1(_01062_),
    .Y(_01076_));
 sky130_fd_sc_hd__a211o_1 _10282_ (.A1(_00929_),
    .A2(_01026_),
    .B1(_01044_),
    .C1(_01057_),
    .X(_01077_));
 sky130_fd_sc_hd__and4_2 _10283_ (.A(_01059_),
    .B(_01075_),
    .C(_01076_),
    .D(_01077_),
    .X(_01078_));
 sky130_fd_sc_hd__o211ai_4 _10284_ (.A1(_01058_),
    .A2(_01078_),
    .B1(_00952_),
    .C1(_01025_),
    .Y(_01079_));
 sky130_fd_sc_hd__a21oi_4 _10285_ (.A1(_00971_),
    .A2(_00972_),
    .B1(_00981_),
    .Y(_01080_));
 sky130_fd_sc_hd__a211o_4 _10286_ (.A1(_01061_),
    .A2(_01076_),
    .B1(_01080_),
    .C1(_00982_),
    .X(_01081_));
 sky130_fd_sc_hd__o211ai_4 _10287_ (.A1(_00982_),
    .A2(_01080_),
    .B1(_01076_),
    .C1(_01061_),
    .Y(_01082_));
 sky130_fd_sc_hd__or3_1 _10288_ (.A(_00966_),
    .B(_00968_),
    .C(_00969_),
    .X(_01083_));
 sky130_fd_sc_hd__nand2_2 _10289_ (.A(_00970_),
    .B(_01083_),
    .Y(_01084_));
 sky130_fd_sc_hd__and4_2 _10290_ (.A(net514),
    .B(net521),
    .C(net768),
    .D(net781),
    .X(_01085_));
 sky130_fd_sc_hd__a22oi_2 _10291_ (.A1(net521),
    .A2(net768),
    .B1(net781),
    .B2(net514),
    .Y(_01086_));
 sky130_fd_sc_hd__and4bb_4 _10292_ (.A_N(_01085_),
    .B_N(_01086_),
    .C(net531),
    .D(net757),
    .X(_01087_));
 sky130_fd_sc_hd__nor2_4 _10293_ (.A(_01085_),
    .B(_01087_),
    .Y(_01088_));
 sky130_fd_sc_hd__o2bb2a_1 _10294_ (.A1_N(net574),
    .A2_N(net722),
    .B1(_00966_),
    .B2(_00967_),
    .X(_01089_));
 sky130_fd_sc_hd__nor2_2 _10295_ (.A(_00968_),
    .B(_01089_),
    .Y(_01090_));
 sky130_fd_sc_hd__or3_4 _10296_ (.A(_00968_),
    .B(_01088_),
    .C(_01089_),
    .X(_01091_));
 sky130_fd_sc_hd__and4_1 _10297_ (.A(net543),
    .B(net557),
    .C(net740),
    .D(net748),
    .X(_01092_));
 sky130_fd_sc_hd__a22oi_2 _10298_ (.A1(net557),
    .A2(net740),
    .B1(net748),
    .B2(net543),
    .Y(_01093_));
 sky130_fd_sc_hd__and4bb_2 _10299_ (.A_N(_01092_),
    .B_N(_01093_),
    .C(net574),
    .D(net731),
    .X(_01094_));
 sky130_fd_sc_hd__or2_4 _10300_ (.A(_01092_),
    .B(_01094_),
    .X(_01095_));
 sky130_fd_sc_hd__xnor2_4 _10301_ (.A(_01088_),
    .B(_01090_),
    .Y(_01096_));
 sky130_fd_sc_hd__nand2_2 _10302_ (.A(_01095_),
    .B(_01096_),
    .Y(_01097_));
 sky130_fd_sc_hd__a21oi_4 _10303_ (.A1(_01091_),
    .A2(_01097_),
    .B1(_01084_),
    .Y(_01098_));
 sky130_fd_sc_hd__a21o_1 _10304_ (.A1(_01091_),
    .A2(_01097_),
    .B1(_01084_),
    .X(_01099_));
 sky130_fd_sc_hd__nand3_2 _10305_ (.A(_01084_),
    .B(_01091_),
    .C(_01097_),
    .Y(_01100_));
 sky130_fd_sc_hd__o2bb2a_1 _10306_ (.A1_N(net595),
    .A2_N(net696),
    .B1(_00975_),
    .B2(_00976_),
    .X(_01101_));
 sky130_fd_sc_hd__nor2_4 _10307_ (.A(_00977_),
    .B(_01101_),
    .Y(_01102_));
 sky130_fd_sc_hd__and2_2 _10308_ (.A(net609),
    .B(net713),
    .X(_01103_));
 sky130_fd_sc_hd__and3_1 _10309_ (.A(net587),
    .B(net696),
    .C(_01103_),
    .X(_01104_));
 sky130_fd_sc_hd__a21oi_1 _10310_ (.A1(net587),
    .A2(net713),
    .B1(_00720_),
    .Y(_01105_));
 sky130_fd_sc_hd__and4bb_2 _10311_ (.A_N(_01104_),
    .B_N(_01105_),
    .C(net599),
    .D(net704),
    .X(_01106_));
 sky130_fd_sc_hd__nor2_2 _10312_ (.A(_01104_),
    .B(_01106_),
    .Y(_01107_));
 sky130_fd_sc_hd__and2b_1 _10313_ (.A_N(_01107_),
    .B(_01102_),
    .X(_01108_));
 sky130_fd_sc_hd__xnor2_4 _10314_ (.A(_01102_),
    .B(_01107_),
    .Y(_01109_));
 sky130_fd_sc_hd__and3_4 _10315_ (.A(_01099_),
    .B(_01100_),
    .C(_01109_),
    .X(_01110_));
 sky130_fd_sc_hd__o211ai_4 _10316_ (.A1(_01098_),
    .A2(_01110_),
    .B1(_01081_),
    .C1(_01082_),
    .Y(_01111_));
 sky130_fd_sc_hd__a211o_2 _10317_ (.A1(_01081_),
    .A2(_01082_),
    .B1(_01098_),
    .C1(_01110_),
    .X(_01112_));
 sky130_fd_sc_hd__a211o_2 _10318_ (.A1(_00952_),
    .A2(_01025_),
    .B1(_01058_),
    .C1(_01078_),
    .X(_01113_));
 sky130_fd_sc_hd__nand4_4 _10319_ (.A(_01079_),
    .B(_01111_),
    .C(_01112_),
    .D(_01113_),
    .Y(_01114_));
 sky130_fd_sc_hd__a211oi_4 _10320_ (.A1(_01079_),
    .A2(_01114_),
    .B1(_00987_),
    .C1(_01024_),
    .Y(_01115_));
 sky130_fd_sc_hd__and4_1 _10321_ (.A(net382),
    .B(net391),
    .C(net901),
    .D(net911),
    .X(_01116_));
 sky130_fd_sc_hd__xnor2_4 _10322_ (.A(_00990_),
    .B(_00992_),
    .Y(_01117_));
 sky130_fd_sc_hd__nand2_2 _10323_ (.A(_01116_),
    .B(_01117_),
    .Y(_01118_));
 sky130_fd_sc_hd__or2_1 _10324_ (.A(_01116_),
    .B(_01117_),
    .X(_01119_));
 sky130_fd_sc_hd__and2_2 _10325_ (.A(_01118_),
    .B(_01119_),
    .X(_01120_));
 sky130_fd_sc_hd__nand3_4 _10326_ (.A(net397),
    .B(net885),
    .C(_01120_),
    .Y(_01121_));
 sky130_fd_sc_hd__a21o_1 _10327_ (.A1(net397),
    .A2(net885),
    .B1(_01120_),
    .X(_01122_));
 sky130_fd_sc_hd__and2_1 _10328_ (.A(_01121_),
    .B(_01122_),
    .X(_01123_));
 sky130_fd_sc_hd__and3_4 _10329_ (.A(_01108_),
    .B(_01121_),
    .C(_01122_),
    .X(_01124_));
 sky130_fd_sc_hd__nand2_4 _10330_ (.A(_01081_),
    .B(_01111_),
    .Y(_01125_));
 sky130_fd_sc_hd__xor2_4 _10331_ (.A(_00979_),
    .B(_01000_),
    .X(_01126_));
 sky130_fd_sc_hd__and2b_1 _10332_ (.A_N(_01126_),
    .B(_01125_),
    .X(_01127_));
 sky130_fd_sc_hd__xnor2_4 _10333_ (.A(_01125_),
    .B(_01126_),
    .Y(_01128_));
 sky130_fd_sc_hd__xnor2_4 _10334_ (.A(_01124_),
    .B(_01128_),
    .Y(_01129_));
 sky130_fd_sc_hd__o211a_2 _10335_ (.A1(_00987_),
    .A2(_01024_),
    .B1(_01079_),
    .C1(_01114_),
    .X(_01130_));
 sky130_fd_sc_hd__nor3_4 _10336_ (.A(_01115_),
    .B(_01129_),
    .C(_01130_),
    .Y(_01131_));
 sky130_fd_sc_hd__o211a_1 _10337_ (.A1(_01115_),
    .A2(_01131_),
    .B1(_01009_),
    .C1(_01023_),
    .X(_01132_));
 sky130_fd_sc_hd__a21o_2 _10338_ (.A1(_01124_),
    .A2(_01128_),
    .B1(_01127_),
    .X(_01133_));
 sky130_fd_sc_hd__a211o_1 _10339_ (.A1(_01009_),
    .A2(_01023_),
    .B1(_01115_),
    .C1(_01131_),
    .X(_01134_));
 sky130_fd_sc_hd__and2b_1 _10340_ (.A_N(_01132_),
    .B(_01134_),
    .X(_01135_));
 sky130_fd_sc_hd__a21o_1 _10341_ (.A1(_01133_),
    .A2(_01134_),
    .B1(_01132_),
    .X(_01136_));
 sky130_fd_sc_hd__and3_2 _10342_ (.A(_01014_),
    .B(_01022_),
    .C(_01136_),
    .X(_01137_));
 sky130_fd_sc_hd__a21oi_4 _10343_ (.A1(_01014_),
    .A2(_01022_),
    .B1(_01136_),
    .Y(_01138_));
 sky130_fd_sc_hd__a211oi_4 _10344_ (.A1(_00863_),
    .A2(_00867_),
    .B1(_01137_),
    .C1(_01138_),
    .Y(_01139_));
 sky130_fd_sc_hd__nor2_2 _10345_ (.A(_01137_),
    .B(_01139_),
    .Y(_01140_));
 sky130_fd_sc_hd__nor2_1 _10346_ (.A(_01021_),
    .B(_01140_),
    .Y(_01141_));
 sky130_fd_sc_hd__or2_1 _10347_ (.A(_01021_),
    .B(_01140_),
    .X(_01142_));
 sky130_fd_sc_hd__or3_4 _10348_ (.A(_00888_),
    .B(_00894_),
    .C(_01019_),
    .X(_01143_));
 sky130_fd_sc_hd__and2_1 _10349_ (.A(_01021_),
    .B(_01140_),
    .X(_01144_));
 sky130_fd_sc_hd__nor2_1 _10350_ (.A(_01141_),
    .B(_01144_),
    .Y(_01145_));
 sky130_fd_sc_hd__o211a_2 _10351_ (.A1(_01137_),
    .A2(_01138_),
    .B1(_00863_),
    .C1(_00867_),
    .X(_01146_));
 sky130_fd_sc_hd__xor2_2 _10352_ (.A(_01133_),
    .B(_01135_),
    .X(_01147_));
 sky130_fd_sc_hd__o21a_2 _10353_ (.A1(_01115_),
    .A2(_01130_),
    .B1(_01129_),
    .X(_01148_));
 sky130_fd_sc_hd__a22o_2 _10354_ (.A1(_01111_),
    .A2(_01112_),
    .B1(_01113_),
    .B2(_01079_),
    .X(_01149_));
 sky130_fd_sc_hd__a22o_1 _10355_ (.A1(_01075_),
    .A2(_01076_),
    .B1(_01077_),
    .B2(_01059_),
    .X(_01150_));
 sky130_fd_sc_hd__nand2b_4 _10356_ (.A_N(_01078_),
    .B(_01150_),
    .Y(_01151_));
 sky130_fd_sc_hd__a21oi_4 _10357_ (.A1(_01043_),
    .A2(_01056_),
    .B1(_01055_),
    .Y(_01152_));
 sky130_fd_sc_hd__xnor2_2 _10358_ (.A(_01040_),
    .B(_01041_),
    .Y(_01153_));
 sky130_fd_sc_hd__nand2_4 _10359_ (.A(net447),
    .B(net863),
    .Y(_01154_));
 sky130_fd_sc_hd__and4_2 _10360_ (.A(net430),
    .B(net439),
    .C(net874),
    .D(net882),
    .X(_01155_));
 sky130_fd_sc_hd__a22oi_1 _10361_ (.A1(net439),
    .A2(net874),
    .B1(net882),
    .B2(net430),
    .Y(_01156_));
 sky130_fd_sc_hd__or2_4 _10362_ (.A(_01155_),
    .B(_01156_),
    .X(_01157_));
 sky130_fd_sc_hd__nor2_2 _10363_ (.A(_01154_),
    .B(_01157_),
    .Y(_01158_));
 sky130_fd_sc_hd__xor2_4 _10364_ (.A(_01154_),
    .B(_01157_),
    .X(_01159_));
 sky130_fd_sc_hd__and2b_2 _10365_ (.A_N(_01031_),
    .B(_01032_),
    .X(_01160_));
 sky130_fd_sc_hd__and3_2 _10366_ (.A(net414),
    .B(net904),
    .C(_01030_),
    .X(_01161_));
 sky130_fd_sc_hd__xnor2_4 _10367_ (.A(_01160_),
    .B(_01161_),
    .Y(_01162_));
 sky130_fd_sc_hd__inv_2 _10368_ (.A(_01162_),
    .Y(_01163_));
 sky130_fd_sc_hd__nand2_1 _10369_ (.A(_01159_),
    .B(_01163_),
    .Y(_01164_));
 sky130_fd_sc_hd__or3_2 _10370_ (.A(_01030_),
    .B(_01033_),
    .C(_01160_),
    .X(_01165_));
 sky130_fd_sc_hd__a21o_4 _10371_ (.A1(_01164_),
    .A2(_01165_),
    .B1(_01153_),
    .X(_01166_));
 sky130_fd_sc_hd__xnor2_2 _10372_ (.A(_01050_),
    .B(_01052_),
    .Y(_01167_));
 sky130_fd_sc_hd__o21ai_4 _10373_ (.A1(_01155_),
    .A2(_01158_),
    .B1(_01167_),
    .Y(_01168_));
 sky130_fd_sc_hd__or3_1 _10374_ (.A(_01155_),
    .B(_01158_),
    .C(_01167_),
    .X(_01169_));
 sky130_fd_sc_hd__and2_2 _10375_ (.A(_01168_),
    .B(_01169_),
    .X(_01170_));
 sky130_fd_sc_hd__and4_1 _10376_ (.A(net457),
    .B(net467),
    .C(net843),
    .D(net853),
    .X(_01171_));
 sky130_fd_sc_hd__nand2_4 _10377_ (.A(net475),
    .B(net834),
    .Y(_01172_));
 sky130_fd_sc_hd__a22oi_4 _10378_ (.A1(net467),
    .A2(net844),
    .B1(net853),
    .B2(net457),
    .Y(_01173_));
 sky130_fd_sc_hd__nor2_2 _10379_ (.A(_01171_),
    .B(_01173_),
    .Y(_01174_));
 sky130_fd_sc_hd__o21ba_1 _10380_ (.A1(_01172_),
    .A2(_01173_),
    .B1_N(_01171_),
    .X(_01175_));
 sky130_fd_sc_hd__nand2b_2 _10381_ (.A_N(_01175_),
    .B(_01170_),
    .Y(_01176_));
 sky130_fd_sc_hd__xnor2_2 _10382_ (.A(_01170_),
    .B(_01175_),
    .Y(_01177_));
 sky130_fd_sc_hd__nand3_2 _10383_ (.A(_01153_),
    .B(_01164_),
    .C(_01165_),
    .Y(_01178_));
 sky130_fd_sc_hd__and3_1 _10384_ (.A(_01166_),
    .B(_01177_),
    .C(_01178_),
    .X(_01179_));
 sky130_fd_sc_hd__nand3_2 _10385_ (.A(_01166_),
    .B(_01177_),
    .C(_01178_),
    .Y(_01180_));
 sky130_fd_sc_hd__a211oi_4 _10386_ (.A1(_01166_),
    .A2(_01180_),
    .B1(_01057_),
    .C1(_01152_),
    .Y(_01181_));
 sky130_fd_sc_hd__nor2_1 _10387_ (.A(_01071_),
    .B(_01073_),
    .Y(_01182_));
 sky130_fd_sc_hd__or2_2 _10388_ (.A(_01074_),
    .B(_01182_),
    .X(_01183_));
 sky130_fd_sc_hd__a21o_4 _10389_ (.A1(_01168_),
    .A2(_01176_),
    .B1(_01183_),
    .X(_01184_));
 sky130_fd_sc_hd__nand3_4 _10390_ (.A(_01168_),
    .B(_01176_),
    .C(_01183_),
    .Y(_01185_));
 sky130_fd_sc_hd__xnor2_4 _10391_ (.A(_01066_),
    .B(_01068_),
    .Y(_01186_));
 sky130_fd_sc_hd__and4_2 _10392_ (.A(net489),
    .B(net499),
    .C(net814),
    .D(net825),
    .X(_01187_));
 sky130_fd_sc_hd__a22oi_2 _10393_ (.A1(net496),
    .A2(net814),
    .B1(net825),
    .B2(net486),
    .Y(_01188_));
 sky130_fd_sc_hd__and4bb_2 _10394_ (.A_N(_01187_),
    .B_N(_01188_),
    .C(net506),
    .D(net804),
    .X(_01189_));
 sky130_fd_sc_hd__nor2_4 _10395_ (.A(_01187_),
    .B(_01189_),
    .Y(_01190_));
 sky130_fd_sc_hd__and2b_1 _10396_ (.A_N(_01190_),
    .B(_01186_),
    .X(_01191_));
 sky130_fd_sc_hd__xnor2_4 _10397_ (.A(_01186_),
    .B(_01190_),
    .Y(_01192_));
 sky130_fd_sc_hd__o2bb2a_1 _10398_ (.A1_N(net531),
    .A2_N(net757),
    .B1(_01085_),
    .B2(_01086_),
    .X(_01193_));
 sky130_fd_sc_hd__nor2_4 _10399_ (.A(_01087_),
    .B(_01193_),
    .Y(_01194_));
 sky130_fd_sc_hd__a21o_2 _10400_ (.A1(_01192_),
    .A2(_01194_),
    .B1(_01191_),
    .X(_01195_));
 sky130_fd_sc_hd__and3_2 _10401_ (.A(_01184_),
    .B(_01185_),
    .C(_01195_),
    .X(_01196_));
 sky130_fd_sc_hd__nand3_4 _10402_ (.A(_01184_),
    .B(_01185_),
    .C(_01195_),
    .Y(_01197_));
 sky130_fd_sc_hd__a21oi_2 _10403_ (.A1(_01184_),
    .A2(_01185_),
    .B1(_01195_),
    .Y(_01198_));
 sky130_fd_sc_hd__o211a_2 _10404_ (.A1(_01057_),
    .A2(_01152_),
    .B1(_01166_),
    .C1(_01180_),
    .X(_01199_));
 sky130_fd_sc_hd__or4_4 _10405_ (.A(_01181_),
    .B(_01196_),
    .C(_01198_),
    .D(_01199_),
    .X(_01200_));
 sky130_fd_sc_hd__and2b_4 _10406_ (.A_N(_01181_),
    .B(_01200_),
    .X(_01201_));
 sky130_fd_sc_hd__nor2_2 _10407_ (.A(_01151_),
    .B(_01201_),
    .Y(_01202_));
 sky130_fd_sc_hd__a21oi_4 _10408_ (.A1(_01099_),
    .A2(_01100_),
    .B1(_01109_),
    .Y(_01203_));
 sky130_fd_sc_hd__a211o_4 _10409_ (.A1(_01184_),
    .A2(_01197_),
    .B1(_01203_),
    .C1(_01110_),
    .X(_01204_));
 sky130_fd_sc_hd__o211ai_4 _10410_ (.A1(_01110_),
    .A2(_01203_),
    .B1(_01197_),
    .C1(_01184_),
    .Y(_01205_));
 sky130_fd_sc_hd__xnor2_4 _10411_ (.A(_01095_),
    .B(_01096_),
    .Y(_01206_));
 sky130_fd_sc_hd__and4_2 _10412_ (.A(net513),
    .B(net520),
    .C(net781),
    .D(net791),
    .X(_01207_));
 sky130_fd_sc_hd__a22oi_2 _10413_ (.A1(net520),
    .A2(net781),
    .B1(net791),
    .B2(net513),
    .Y(_01208_));
 sky130_fd_sc_hd__and4bb_2 _10414_ (.A_N(_01207_),
    .B_N(_01208_),
    .C(net529),
    .D(net769),
    .X(_01209_));
 sky130_fd_sc_hd__nor2_4 _10415_ (.A(_01207_),
    .B(_01209_),
    .Y(_01210_));
 sky130_fd_sc_hd__o2bb2a_1 _10416_ (.A1_N(net574),
    .A2_N(net731),
    .B1(_01092_),
    .B2(_01093_),
    .X(_01211_));
 sky130_fd_sc_hd__nor2_2 _10417_ (.A(_01094_),
    .B(_01211_),
    .Y(_01212_));
 sky130_fd_sc_hd__or3_4 _10418_ (.A(_01094_),
    .B(_01210_),
    .C(_01211_),
    .X(_01213_));
 sky130_fd_sc_hd__and4_1 _10419_ (.A(net541),
    .B(net555),
    .C(net748),
    .D(net757),
    .X(_01214_));
 sky130_fd_sc_hd__a22oi_2 _10420_ (.A1(net555),
    .A2(net748),
    .B1(net757),
    .B2(net541),
    .Y(_01215_));
 sky130_fd_sc_hd__and4bb_2 _10421_ (.A_N(_01214_),
    .B_N(_01215_),
    .C(net572),
    .D(net740),
    .X(_01216_));
 sky130_fd_sc_hd__or2_4 _10422_ (.A(_01214_),
    .B(_01216_),
    .X(_01217_));
 sky130_fd_sc_hd__xnor2_4 _10423_ (.A(_01210_),
    .B(_01212_),
    .Y(_01218_));
 sky130_fd_sc_hd__nand2_2 _10424_ (.A(_01217_),
    .B(_01218_),
    .Y(_01219_));
 sky130_fd_sc_hd__a21oi_4 _10425_ (.A1(_01213_),
    .A2(_01219_),
    .B1(_01206_),
    .Y(_01220_));
 sky130_fd_sc_hd__a21o_1 _10426_ (.A1(_01213_),
    .A2(_01219_),
    .B1(_01206_),
    .X(_01221_));
 sky130_fd_sc_hd__nand3_2 _10427_ (.A(_01206_),
    .B(_01213_),
    .C(_01219_),
    .Y(_01222_));
 sky130_fd_sc_hd__o2bb2a_1 _10428_ (.A1_N(net599),
    .A2_N(net705),
    .B1(_01104_),
    .B2(_01105_),
    .X(_01223_));
 sky130_fd_sc_hd__nor2_4 _10429_ (.A(_01106_),
    .B(_01223_),
    .Y(_01224_));
 sky130_fd_sc_hd__and2_2 _10430_ (.A(net609),
    .B(net722),
    .X(_01225_));
 sky130_fd_sc_hd__and3_2 _10431_ (.A(net587),
    .B(net705),
    .C(_01225_),
    .X(_01226_));
 sky130_fd_sc_hd__a21oi_1 _10432_ (.A1(net581),
    .A2(net722),
    .B1(_00974_),
    .Y(_01227_));
 sky130_fd_sc_hd__and4bb_2 _10433_ (.A_N(_01226_),
    .B_N(_01227_),
    .C(net599),
    .D(net713),
    .X(_01228_));
 sky130_fd_sc_hd__nor2_4 _10434_ (.A(_01226_),
    .B(_01228_),
    .Y(_01229_));
 sky130_fd_sc_hd__and2b_1 _10435_ (.A_N(_01229_),
    .B(_01224_),
    .X(_01230_));
 sky130_fd_sc_hd__xnor2_4 _10436_ (.A(_01224_),
    .B(_01229_),
    .Y(_01231_));
 sky130_fd_sc_hd__and3_4 _10437_ (.A(_01221_),
    .B(_01222_),
    .C(_01231_),
    .X(_01232_));
 sky130_fd_sc_hd__a211o_1 _10438_ (.A1(_01204_),
    .A2(_01205_),
    .B1(_01220_),
    .C1(_01232_),
    .X(_01233_));
 sky130_fd_sc_hd__o211ai_4 _10439_ (.A1(_01220_),
    .A2(_01232_),
    .B1(_01204_),
    .C1(_01205_),
    .Y(_01234_));
 sky130_fd_sc_hd__nand2_4 _10440_ (.A(_01233_),
    .B(_01234_),
    .Y(_01235_));
 sky130_fd_sc_hd__xnor2_4 _10441_ (.A(_01151_),
    .B(_01201_),
    .Y(_01236_));
 sky130_fd_sc_hd__nor2_2 _10442_ (.A(_01235_),
    .B(_01236_),
    .Y(_01237_));
 sky130_fd_sc_hd__o211ai_4 _10443_ (.A1(_01202_),
    .A2(_01237_),
    .B1(_01114_),
    .C1(_01149_),
    .Y(_01238_));
 sky130_fd_sc_hd__a22oi_1 _10444_ (.A1(net391),
    .A2(net904),
    .B1(net910),
    .B2(net382),
    .Y(_01239_));
 sky130_fd_sc_hd__nor2_1 _10445_ (.A(_01116_),
    .B(_01239_),
    .Y(_01240_));
 sky130_fd_sc_hd__and3_2 _10446_ (.A(net397),
    .B(net896),
    .C(_01240_),
    .X(_01241_));
 sky130_fd_sc_hd__a21oi_1 _10447_ (.A1(net397),
    .A2(net896),
    .B1(_01240_),
    .Y(_01242_));
 sky130_fd_sc_hd__nor2_2 _10448_ (.A(_01241_),
    .B(_01242_),
    .Y(_01243_));
 sky130_fd_sc_hd__nand2_4 _10449_ (.A(_01230_),
    .B(_01243_),
    .Y(_01244_));
 sky130_fd_sc_hd__nor2_1 _10450_ (.A(_01108_),
    .B(_01123_),
    .Y(_01245_));
 sky130_fd_sc_hd__or2_1 _10451_ (.A(_01124_),
    .B(_01245_),
    .X(_01246_));
 sky130_fd_sc_hd__a21o_2 _10452_ (.A1(_01204_),
    .A2(_01234_),
    .B1(_01246_),
    .X(_01247_));
 sky130_fd_sc_hd__nand3_1 _10453_ (.A(_01204_),
    .B(_01234_),
    .C(_01246_),
    .Y(_01248_));
 sky130_fd_sc_hd__nand2_2 _10454_ (.A(_01247_),
    .B(_01248_),
    .Y(_01249_));
 sky130_fd_sc_hd__or2_2 _10455_ (.A(_01244_),
    .B(_01249_),
    .X(_01250_));
 sky130_fd_sc_hd__xor2_4 _10456_ (.A(_01244_),
    .B(_01249_),
    .X(_01251_));
 sky130_fd_sc_hd__a211o_4 _10457_ (.A1(_01114_),
    .A2(_01149_),
    .B1(_01202_),
    .C1(_01237_),
    .X(_01252_));
 sky130_fd_sc_hd__and3_2 _10458_ (.A(_01238_),
    .B(_01251_),
    .C(_01252_),
    .X(_01253_));
 sky130_fd_sc_hd__nand3_4 _10459_ (.A(_01238_),
    .B(_01251_),
    .C(_01252_),
    .Y(_01254_));
 sky130_fd_sc_hd__a211oi_4 _10460_ (.A1(_01238_),
    .A2(_01254_),
    .B1(_01131_),
    .C1(_01148_),
    .Y(_01255_));
 sky130_fd_sc_hd__o211a_2 _10461_ (.A1(_01131_),
    .A2(_01148_),
    .B1(_01238_),
    .C1(_01254_),
    .X(_01256_));
 sky130_fd_sc_hd__a211oi_4 _10462_ (.A1(_01247_),
    .A2(_01250_),
    .B1(_01255_),
    .C1(_01256_),
    .Y(_01257_));
 sky130_fd_sc_hd__nor2_2 _10463_ (.A(_01255_),
    .B(_01257_),
    .Y(_01258_));
 sky130_fd_sc_hd__and2b_1 _10464_ (.A_N(_01258_),
    .B(_01147_),
    .X(_01259_));
 sky130_fd_sc_hd__xnor2_1 _10465_ (.A(_01147_),
    .B(_01258_),
    .Y(_01260_));
 sky130_fd_sc_hd__o21a_1 _10466_ (.A1(_00996_),
    .A2(_00998_),
    .B1(_01260_),
    .X(_01261_));
 sky130_fd_sc_hd__nor2_2 _10467_ (.A(_01259_),
    .B(_01261_),
    .Y(_01262_));
 sky130_fd_sc_hd__o21ai_4 _10468_ (.A1(_01139_),
    .A2(_01146_),
    .B1(_01262_),
    .Y(_01263_));
 sky130_fd_sc_hd__nor3_1 _10469_ (.A(_00996_),
    .B(_00998_),
    .C(_01260_),
    .Y(_01264_));
 sky130_fd_sc_hd__or2_2 _10470_ (.A(_01261_),
    .B(_01264_),
    .X(_01265_));
 sky130_fd_sc_hd__o211a_2 _10471_ (.A1(_01255_),
    .A2(_01256_),
    .B1(_01247_),
    .C1(_01250_),
    .X(_01266_));
 sky130_fd_sc_hd__a21oi_4 _10472_ (.A1(_01238_),
    .A2(_01252_),
    .B1(_01251_),
    .Y(_01267_));
 sky130_fd_sc_hd__xnor2_4 _10473_ (.A(_01235_),
    .B(_01236_),
    .Y(_01268_));
 sky130_fd_sc_hd__o22ai_4 _10474_ (.A1(_01196_),
    .A2(_01198_),
    .B1(_01199_),
    .B2(_01181_),
    .Y(_01269_));
 sky130_fd_sc_hd__a21oi_2 _10475_ (.A1(_01166_),
    .A2(_01178_),
    .B1(_01177_),
    .Y(_01270_));
 sky130_fd_sc_hd__a22oi_4 _10476_ (.A1(net440),
    .A2(net883),
    .B1(net894),
    .B2(net431),
    .Y(_01271_));
 sky130_fd_sc_hd__and4_1 _10477_ (.A(net431),
    .B(net440),
    .C(net883),
    .D(net894),
    .X(_01272_));
 sky130_fd_sc_hd__nor2_2 _10478_ (.A(_01271_),
    .B(_01272_),
    .Y(_01273_));
 sky130_fd_sc_hd__nand2_2 _10479_ (.A(net447),
    .B(net873),
    .Y(_01274_));
 sky130_fd_sc_hd__xnor2_4 _10480_ (.A(_01273_),
    .B(_01274_),
    .Y(_01275_));
 sky130_fd_sc_hd__a22o_1 _10481_ (.A1(net422),
    .A2(net904),
    .B1(net913),
    .B2(net414),
    .X(_01276_));
 sky130_fd_sc_hd__o21a_2 _10482_ (.A1(_01030_),
    .A2(_01033_),
    .B1(_01276_),
    .X(_01277_));
 sky130_fd_sc_hd__nand2_1 _10483_ (.A(_01275_),
    .B(_01277_),
    .Y(_01278_));
 sky130_fd_sc_hd__xor2_2 _10484_ (.A(_01159_),
    .B(_01162_),
    .X(_01279_));
 sky130_fd_sc_hd__or2_1 _10485_ (.A(_01278_),
    .B(_01279_),
    .X(_01280_));
 sky130_fd_sc_hd__o21ba_2 _10486_ (.A1(_01271_),
    .A2(_01274_),
    .B1_N(_01272_),
    .X(_01281_));
 sky130_fd_sc_hd__xnor2_4 _10487_ (.A(_01172_),
    .B(_01174_),
    .Y(_01282_));
 sky130_fd_sc_hd__nand2b_2 _10488_ (.A_N(_01281_),
    .B(_01282_),
    .Y(_01283_));
 sky130_fd_sc_hd__xnor2_2 _10489_ (.A(_01281_),
    .B(_01282_),
    .Y(_01284_));
 sky130_fd_sc_hd__and4_1 _10490_ (.A(net456),
    .B(net466),
    .C(net853),
    .D(net864),
    .X(_01285_));
 sky130_fd_sc_hd__nand2_4 _10491_ (.A(net475),
    .B(net844),
    .Y(_01286_));
 sky130_fd_sc_hd__a22oi_4 _10492_ (.A1(net466),
    .A2(net853),
    .B1(net869),
    .B2(net456),
    .Y(_01287_));
 sky130_fd_sc_hd__nor2_2 _10493_ (.A(_01285_),
    .B(_01287_),
    .Y(_01288_));
 sky130_fd_sc_hd__o21ba_1 _10494_ (.A1(_01286_),
    .A2(_01287_),
    .B1_N(_01285_),
    .X(_01289_));
 sky130_fd_sc_hd__nand2b_2 _10495_ (.A_N(_01289_),
    .B(_01284_),
    .Y(_01290_));
 sky130_fd_sc_hd__xor2_1 _10496_ (.A(_01284_),
    .B(_01289_),
    .X(_01291_));
 sky130_fd_sc_hd__xnor2_1 _10497_ (.A(_01278_),
    .B(_01279_),
    .Y(_01292_));
 sky130_fd_sc_hd__or2_2 _10498_ (.A(_01291_),
    .B(_01292_),
    .X(_01293_));
 sky130_fd_sc_hd__clkinv_2 _10499_ (.A(_01293_),
    .Y(_01294_));
 sky130_fd_sc_hd__a211oi_2 _10500_ (.A1(_01280_),
    .A2(_01293_),
    .B1(_01179_),
    .C1(_01270_),
    .Y(_01295_));
 sky130_fd_sc_hd__xnor2_4 _10501_ (.A(_01192_),
    .B(_01194_),
    .Y(_01296_));
 sky130_fd_sc_hd__a21o_4 _10502_ (.A1(_01283_),
    .A2(_01290_),
    .B1(_01296_),
    .X(_01297_));
 sky130_fd_sc_hd__nand3_2 _10503_ (.A(_01283_),
    .B(_01290_),
    .C(_01296_),
    .Y(_01298_));
 sky130_fd_sc_hd__o2bb2a_1 _10504_ (.A1_N(net506),
    .A2_N(net804),
    .B1(_01187_),
    .B2(_01188_),
    .X(_01299_));
 sky130_fd_sc_hd__nor2_2 _10505_ (.A(_01189_),
    .B(_01299_),
    .Y(_01300_));
 sky130_fd_sc_hd__and4_1 _10506_ (.A(net486),
    .B(net496),
    .C(net825),
    .D(net834),
    .X(_01301_));
 sky130_fd_sc_hd__a22oi_2 _10507_ (.A1(net496),
    .A2(net825),
    .B1(net834),
    .B2(net486),
    .Y(_01302_));
 sky130_fd_sc_hd__and4bb_2 _10508_ (.A_N(_01301_),
    .B_N(_01302_),
    .C(net504),
    .D(net814),
    .X(_01303_));
 sky130_fd_sc_hd__nor2_2 _10509_ (.A(_01301_),
    .B(_01303_),
    .Y(_01304_));
 sky130_fd_sc_hd__and2b_2 _10510_ (.A_N(_01304_),
    .B(_01300_),
    .X(_01305_));
 sky130_fd_sc_hd__xnor2_2 _10511_ (.A(_01300_),
    .B(_01304_),
    .Y(_01306_));
 sky130_fd_sc_hd__o2bb2a_1 _10512_ (.A1_N(net529),
    .A2_N(net769),
    .B1(_01207_),
    .B2(_01208_),
    .X(_01307_));
 sky130_fd_sc_hd__nor2_2 _10513_ (.A(_01209_),
    .B(_01307_),
    .Y(_01308_));
 sky130_fd_sc_hd__and2_2 _10514_ (.A(_01306_),
    .B(_01308_),
    .X(_01309_));
 sky130_fd_sc_hd__o211ai_4 _10515_ (.A1(_01305_),
    .A2(_01309_),
    .B1(_01297_),
    .C1(_01298_),
    .Y(_01310_));
 sky130_fd_sc_hd__a211o_1 _10516_ (.A1(_01297_),
    .A2(_01298_),
    .B1(_01305_),
    .C1(_01309_),
    .X(_01311_));
 sky130_fd_sc_hd__nand2_2 _10517_ (.A(_01310_),
    .B(_01311_),
    .Y(_01312_));
 sky130_fd_sc_hd__o211a_2 _10518_ (.A1(_01179_),
    .A2(_01270_),
    .B1(_01280_),
    .C1(_01293_),
    .X(_01313_));
 sky130_fd_sc_hd__nor3_4 _10519_ (.A(net122),
    .B(_01312_),
    .C(_01313_),
    .Y(_01314_));
 sky130_fd_sc_hd__o211a_4 _10520_ (.A1(net122),
    .A2(_01314_),
    .B1(_01200_),
    .C1(_01269_),
    .X(_01315_));
 sky130_fd_sc_hd__a21oi_4 _10521_ (.A1(_01221_),
    .A2(_01222_),
    .B1(_01231_),
    .Y(_01316_));
 sky130_fd_sc_hd__a211o_4 _10522_ (.A1(_01297_),
    .A2(_01310_),
    .B1(_01316_),
    .C1(_01232_),
    .X(_01317_));
 sky130_fd_sc_hd__o211ai_4 _10523_ (.A1(_01232_),
    .A2(_01316_),
    .B1(_01310_),
    .C1(_01297_),
    .Y(_01318_));
 sky130_fd_sc_hd__xnor2_4 _10524_ (.A(_01217_),
    .B(_01218_),
    .Y(_01319_));
 sky130_fd_sc_hd__and4_2 _10525_ (.A(net513),
    .B(net520),
    .C(net791),
    .D(net804),
    .X(_01320_));
 sky130_fd_sc_hd__a22oi_2 _10526_ (.A1(net520),
    .A2(net791),
    .B1(net804),
    .B2(net513),
    .Y(_01321_));
 sky130_fd_sc_hd__and4bb_2 _10527_ (.A_N(_01320_),
    .B_N(_01321_),
    .C(net529),
    .D(net781),
    .X(_01322_));
 sky130_fd_sc_hd__nor2_4 _10528_ (.A(_01320_),
    .B(_01322_),
    .Y(_01323_));
 sky130_fd_sc_hd__o2bb2a_1 _10529_ (.A1_N(net572),
    .A2_N(net740),
    .B1(_01214_),
    .B2(_01215_),
    .X(_01324_));
 sky130_fd_sc_hd__nor2_2 _10530_ (.A(_01216_),
    .B(_01324_),
    .Y(_01325_));
 sky130_fd_sc_hd__or3_4 _10531_ (.A(_01216_),
    .B(_01323_),
    .C(_01324_),
    .X(_01326_));
 sky130_fd_sc_hd__and4_1 _10532_ (.A(net541),
    .B(net555),
    .C(net757),
    .D(net768),
    .X(_01327_));
 sky130_fd_sc_hd__a22oi_2 _10533_ (.A1(net555),
    .A2(net757),
    .B1(net768),
    .B2(net541),
    .Y(_01328_));
 sky130_fd_sc_hd__and4bb_2 _10534_ (.A_N(_01327_),
    .B_N(_01328_),
    .C(net572),
    .D(net748),
    .X(_01329_));
 sky130_fd_sc_hd__or2_4 _10535_ (.A(_01327_),
    .B(_01329_),
    .X(_01330_));
 sky130_fd_sc_hd__xnor2_4 _10536_ (.A(_01323_),
    .B(_01325_),
    .Y(_01331_));
 sky130_fd_sc_hd__nand2_2 _10537_ (.A(_01330_),
    .B(_01331_),
    .Y(_01332_));
 sky130_fd_sc_hd__a21oi_4 _10538_ (.A1(_01326_),
    .A2(_01332_),
    .B1(_01319_),
    .Y(_01333_));
 sky130_fd_sc_hd__a21o_1 _10539_ (.A1(_01326_),
    .A2(_01332_),
    .B1(_01319_),
    .X(_01334_));
 sky130_fd_sc_hd__nand3_2 _10540_ (.A(_01319_),
    .B(_01326_),
    .C(_01332_),
    .Y(_01335_));
 sky130_fd_sc_hd__o2bb2a_1 _10541_ (.A1_N(net599),
    .A2_N(net714),
    .B1(_01226_),
    .B2(_01227_),
    .X(_01336_));
 sky130_fd_sc_hd__and2_4 _10542_ (.A(net615),
    .B(net732),
    .X(_01337_));
 sky130_fd_sc_hd__and3_1 _10543_ (.A(net587),
    .B(net714),
    .C(_01337_),
    .X(_01338_));
 sky130_fd_sc_hd__a21oi_1 _10544_ (.A1(net587),
    .A2(net731),
    .B1(_01103_),
    .Y(_01339_));
 sky130_fd_sc_hd__and4bb_2 _10545_ (.A_N(_01338_),
    .B_N(_01339_),
    .C(net599),
    .D(net722),
    .X(_01340_));
 sky130_fd_sc_hd__nor2_1 _10546_ (.A(_01338_),
    .B(_01340_),
    .Y(_01341_));
 sky130_fd_sc_hd__or3_1 _10547_ (.A(_01228_),
    .B(_01336_),
    .C(_01341_),
    .X(_01342_));
 sky130_fd_sc_hd__o21ai_1 _10548_ (.A1(_01228_),
    .A2(_01336_),
    .B1(_01341_),
    .Y(_01343_));
 sky130_fd_sc_hd__and2_2 _10549_ (.A(_01342_),
    .B(_01343_),
    .X(_01344_));
 sky130_fd_sc_hd__and3_4 _10550_ (.A(_01334_),
    .B(_01335_),
    .C(_01344_),
    .X(_01345_));
 sky130_fd_sc_hd__o211ai_4 _10551_ (.A1(_01333_),
    .A2(_01345_),
    .B1(_01317_),
    .C1(_01318_),
    .Y(_01346_));
 sky130_fd_sc_hd__a211o_1 _10552_ (.A1(_01317_),
    .A2(_01318_),
    .B1(_01333_),
    .C1(_01345_),
    .X(_01347_));
 sky130_fd_sc_hd__nand2_2 _10553_ (.A(_01346_),
    .B(_01347_),
    .Y(_01348_));
 sky130_fd_sc_hd__a211oi_4 _10554_ (.A1(_01200_),
    .A2(_01269_),
    .B1(net122),
    .C1(_01314_),
    .Y(_01349_));
 sky130_fd_sc_hd__or3_4 _10555_ (.A(_01315_),
    .B(_01348_),
    .C(_01349_),
    .X(_01350_));
 sky130_fd_sc_hd__and2b_2 _10556_ (.A_N(_01315_),
    .B(_01350_),
    .X(_01351_));
 sky130_fd_sc_hd__or2_2 _10557_ (.A(_01268_),
    .B(_01351_),
    .X(_01352_));
 sky130_fd_sc_hd__a22oi_1 _10558_ (.A1(net398),
    .A2(net909),
    .B1(net915),
    .B2(net391),
    .Y(_01353_));
 sky130_fd_sc_hd__nand2_1 _10559_ (.A(net398),
    .B(net915),
    .Y(_01354_));
 sky130_fd_sc_hd__and4_4 _10560_ (.A(net391),
    .B(net398),
    .C(net909),
    .D(net915),
    .X(_01355_));
 sky130_fd_sc_hd__or2_1 _10561_ (.A(_01353_),
    .B(_01355_),
    .X(_01356_));
 sky130_fd_sc_hd__or2_2 _10562_ (.A(_01342_),
    .B(_01356_),
    .X(_01357_));
 sky130_fd_sc_hd__or2_1 _10563_ (.A(_01230_),
    .B(_01243_),
    .X(_01358_));
 sky130_fd_sc_hd__nand2_2 _10564_ (.A(_01244_),
    .B(_01358_),
    .Y(_01359_));
 sky130_fd_sc_hd__a21oi_4 _10565_ (.A1(_01317_),
    .A2(_01346_),
    .B1(_01359_),
    .Y(_01360_));
 sky130_fd_sc_hd__and3_1 _10566_ (.A(_01317_),
    .B(_01346_),
    .C(_01359_),
    .X(_01361_));
 sky130_fd_sc_hd__or2_2 _10567_ (.A(_01360_),
    .B(_01361_),
    .X(_01362_));
 sky130_fd_sc_hd__nor2_4 _10568_ (.A(_01357_),
    .B(_01362_),
    .Y(_01363_));
 sky130_fd_sc_hd__and2_1 _10569_ (.A(_01357_),
    .B(_01362_),
    .X(_01364_));
 sky130_fd_sc_hd__nor2_2 _10570_ (.A(_01363_),
    .B(_01364_),
    .Y(_01365_));
 sky130_fd_sc_hd__xnor2_4 _10571_ (.A(_01268_),
    .B(_01351_),
    .Y(_01366_));
 sky130_fd_sc_hd__or3_4 _10572_ (.A(_01363_),
    .B(_01364_),
    .C(_01366_),
    .X(_01367_));
 sky130_fd_sc_hd__a211o_4 _10573_ (.A1(_01352_),
    .A2(_01367_),
    .B1(_01253_),
    .C1(_01267_),
    .X(_01368_));
 sky130_fd_sc_hd__o211ai_4 _10574_ (.A1(_01253_),
    .A2(_01267_),
    .B1(_01352_),
    .C1(_01367_),
    .Y(_01369_));
 sky130_fd_sc_hd__o211ai_4 _10575_ (.A1(_01360_),
    .A2(_01363_),
    .B1(_01368_),
    .C1(_01369_),
    .Y(_01370_));
 sky130_fd_sc_hd__a211oi_4 _10576_ (.A1(_01368_),
    .A2(_01370_),
    .B1(_01257_),
    .C1(_01266_),
    .Y(_01371_));
 sky130_fd_sc_hd__o211a_2 _10577_ (.A1(_01257_),
    .A2(_01266_),
    .B1(_01368_),
    .C1(_01370_),
    .X(_01372_));
 sky130_fd_sc_hd__a211oi_4 _10578_ (.A1(_01118_),
    .A2(_01121_),
    .B1(_01371_),
    .C1(_01372_),
    .Y(_01373_));
 sky130_fd_sc_hd__nor2_1 _10579_ (.A(_01371_),
    .B(_01373_),
    .Y(_01374_));
 sky130_fd_sc_hd__or2_1 _10580_ (.A(_01265_),
    .B(_01374_),
    .X(_01375_));
 sky130_fd_sc_hd__or3_4 _10581_ (.A(_01139_),
    .B(_01146_),
    .C(_01262_),
    .X(_01376_));
 sky130_fd_sc_hd__nand2_1 _10582_ (.A(_01265_),
    .B(_01374_),
    .Y(_01377_));
 sky130_fd_sc_hd__and2_4 _10583_ (.A(_01375_),
    .B(_01377_),
    .X(_01378_));
 sky130_fd_sc_hd__o211a_1 _10584_ (.A1(_01371_),
    .A2(_01372_),
    .B1(_01118_),
    .C1(_01121_),
    .X(_01379_));
 sky130_fd_sc_hd__a211o_2 _10585_ (.A1(_01368_),
    .A2(_01369_),
    .B1(_01360_),
    .C1(_01363_),
    .X(_01380_));
 sky130_fd_sc_hd__xnor2_4 _10586_ (.A(_01365_),
    .B(_01366_),
    .Y(_01381_));
 sky130_fd_sc_hd__o21ai_4 _10587_ (.A1(_01315_),
    .A2(_01349_),
    .B1(_01348_),
    .Y(_01382_));
 sky130_fd_sc_hd__o21a_1 _10588_ (.A1(_01295_),
    .A2(_01313_),
    .B1(_01312_),
    .X(_01383_));
 sky130_fd_sc_hd__and2_2 _10589_ (.A(_01291_),
    .B(_01292_),
    .X(_01384_));
 sky130_fd_sc_hd__a22o_1 _10590_ (.A1(net440),
    .A2(net895),
    .B1(net903),
    .B2(net430),
    .X(_01385_));
 sky130_fd_sc_hd__and4_1 _10591_ (.A(net430),
    .B(net440),
    .C(net895),
    .D(net903),
    .X(_01386_));
 sky130_fd_sc_hd__inv_2 _10592_ (.A(_01386_),
    .Y(_01387_));
 sky130_fd_sc_hd__nand2_2 _10593_ (.A(_01385_),
    .B(_01387_),
    .Y(_01388_));
 sky130_fd_sc_hd__nand2_2 _10594_ (.A(net447),
    .B(net883),
    .Y(_01389_));
 sky130_fd_sc_hd__xnor2_4 _10595_ (.A(_01388_),
    .B(_01389_),
    .Y(_01390_));
 sky130_fd_sc_hd__or2_4 _10596_ (.A(_01030_),
    .B(_01390_),
    .X(_01391_));
 sky130_fd_sc_hd__xnor2_4 _10597_ (.A(_01275_),
    .B(_01277_),
    .Y(_01392_));
 sky130_fd_sc_hd__or2_2 _10598_ (.A(_01391_),
    .B(_01392_),
    .X(_01393_));
 sky130_fd_sc_hd__xor2_4 _10599_ (.A(_01391_),
    .B(_01392_),
    .X(_01394_));
 sky130_fd_sc_hd__a31o_4 _10600_ (.A1(net447),
    .A2(net883),
    .A3(_01385_),
    .B1(_01386_),
    .X(_01395_));
 sky130_fd_sc_hd__xnor2_4 _10601_ (.A(_01286_),
    .B(_01288_),
    .Y(_01396_));
 sky130_fd_sc_hd__nand2_1 _10602_ (.A(_01395_),
    .B(_01396_),
    .Y(_01397_));
 sky130_fd_sc_hd__xor2_4 _10603_ (.A(_01395_),
    .B(_01396_),
    .X(_01398_));
 sky130_fd_sc_hd__and4_1 _10604_ (.A(net456),
    .B(net466),
    .C(net869),
    .D(net873),
    .X(_01399_));
 sky130_fd_sc_hd__nand2_4 _10605_ (.A(net475),
    .B(net853),
    .Y(_01400_));
 sky130_fd_sc_hd__a22oi_4 _10606_ (.A1(net466),
    .A2(net864),
    .B1(net873),
    .B2(net456),
    .Y(_01401_));
 sky130_fd_sc_hd__nor2_2 _10607_ (.A(_01399_),
    .B(_01401_),
    .Y(_01402_));
 sky130_fd_sc_hd__o21ba_2 _10608_ (.A1(_01400_),
    .A2(_01401_),
    .B1_N(_01399_),
    .X(_01403_));
 sky130_fd_sc_hd__nand2b_2 _10609_ (.A_N(_01403_),
    .B(_01398_),
    .Y(_01404_));
 sky130_fd_sc_hd__xnor2_4 _10610_ (.A(_01398_),
    .B(_01403_),
    .Y(_01405_));
 sky130_fd_sc_hd__nand2_2 _10611_ (.A(_01394_),
    .B(_01405_),
    .Y(_01406_));
 sky130_fd_sc_hd__a211o_4 _10612_ (.A1(_01393_),
    .A2(_01406_),
    .B1(_01294_),
    .C1(_01384_),
    .X(_01407_));
 sky130_fd_sc_hd__xnor2_2 _10613_ (.A(_01306_),
    .B(_01308_),
    .Y(_01408_));
 sky130_fd_sc_hd__a21o_4 _10614_ (.A1(_01397_),
    .A2(_01404_),
    .B1(_01408_),
    .X(_01409_));
 sky130_fd_sc_hd__nand3_2 _10615_ (.A(_01397_),
    .B(_01404_),
    .C(_01408_),
    .Y(_01410_));
 sky130_fd_sc_hd__o2bb2a_1 _10616_ (.A1_N(net504),
    .A2_N(net814),
    .B1(_01301_),
    .B2(_01302_),
    .X(_01411_));
 sky130_fd_sc_hd__nor2_2 _10617_ (.A(_01303_),
    .B(_01411_),
    .Y(_01412_));
 sky130_fd_sc_hd__and4_1 _10618_ (.A(net486),
    .B(net496),
    .C(net833),
    .D(net843),
    .X(_01413_));
 sky130_fd_sc_hd__nand2_8 _10619_ (.A(net505),
    .B(net827),
    .Y(_01414_));
 sky130_fd_sc_hd__a22oi_4 _10620_ (.A1(net496),
    .A2(net833),
    .B1(net843),
    .B2(net486),
    .Y(_01415_));
 sky130_fd_sc_hd__nor2_2 _10621_ (.A(_01413_),
    .B(_01415_),
    .Y(_01416_));
 sky130_fd_sc_hd__o21ba_1 _10622_ (.A1(_01414_),
    .A2(_01415_),
    .B1_N(_01413_),
    .X(_01417_));
 sky130_fd_sc_hd__and2b_2 _10623_ (.A_N(_01417_),
    .B(_01412_),
    .X(_01418_));
 sky130_fd_sc_hd__xnor2_2 _10624_ (.A(_01412_),
    .B(_01417_),
    .Y(_01419_));
 sky130_fd_sc_hd__o2bb2a_1 _10625_ (.A1_N(net529),
    .A2_N(net781),
    .B1(_01320_),
    .B2(_01321_),
    .X(_01420_));
 sky130_fd_sc_hd__nor2_2 _10626_ (.A(_01322_),
    .B(_01420_),
    .Y(_01421_));
 sky130_fd_sc_hd__and2_2 _10627_ (.A(_01419_),
    .B(_01421_),
    .X(_01422_));
 sky130_fd_sc_hd__o211ai_4 _10628_ (.A1(_01418_),
    .A2(_01422_),
    .B1(_01409_),
    .C1(_01410_),
    .Y(_01423_));
 sky130_fd_sc_hd__a211o_2 _10629_ (.A1(_01409_),
    .A2(_01410_),
    .B1(_01418_),
    .C1(_01422_),
    .X(_01424_));
 sky130_fd_sc_hd__o211ai_4 _10630_ (.A1(_01294_),
    .A2(_01384_),
    .B1(_01393_),
    .C1(_01406_),
    .Y(_01425_));
 sky130_fd_sc_hd__and4_2 _10631_ (.A(_01407_),
    .B(_01423_),
    .C(_01424_),
    .D(_01425_),
    .X(_01426_));
 sky130_fd_sc_hd__nand4_2 _10632_ (.A(_01407_),
    .B(_01423_),
    .C(_01424_),
    .D(_01425_),
    .Y(_01427_));
 sky130_fd_sc_hd__a211oi_2 _10633_ (.A1(_01407_),
    .A2(_01427_),
    .B1(_01314_),
    .C1(_01383_),
    .Y(_01428_));
 sky130_fd_sc_hd__a21oi_4 _10634_ (.A1(_01334_),
    .A2(_01335_),
    .B1(_01344_),
    .Y(_01429_));
 sky130_fd_sc_hd__a211o_4 _10635_ (.A1(_01409_),
    .A2(_01423_),
    .B1(_01429_),
    .C1(_01345_),
    .X(_01430_));
 sky130_fd_sc_hd__o211ai_4 _10636_ (.A1(_01345_),
    .A2(_01429_),
    .B1(_01423_),
    .C1(_01409_),
    .Y(_01431_));
 sky130_fd_sc_hd__xnor2_4 _10637_ (.A(_01330_),
    .B(_01331_),
    .Y(_01432_));
 sky130_fd_sc_hd__and4_2 _10638_ (.A(net513),
    .B(net520),
    .C(net804),
    .D(net814),
    .X(_01433_));
 sky130_fd_sc_hd__a22oi_2 _10639_ (.A1(net520),
    .A2(net804),
    .B1(net814),
    .B2(net513),
    .Y(_01434_));
 sky130_fd_sc_hd__and4bb_4 _10640_ (.A_N(_01433_),
    .B_N(_01434_),
    .C(net529),
    .D(net791),
    .X(_01435_));
 sky130_fd_sc_hd__nor2_4 _10641_ (.A(_01433_),
    .B(_01435_),
    .Y(_01436_));
 sky130_fd_sc_hd__o2bb2a_1 _10642_ (.A1_N(net572),
    .A2_N(net748),
    .B1(_01327_),
    .B2(_01328_),
    .X(_01437_));
 sky130_fd_sc_hd__nor2_2 _10643_ (.A(_01329_),
    .B(_01437_),
    .Y(_01438_));
 sky130_fd_sc_hd__or3_4 _10644_ (.A(_01329_),
    .B(_01436_),
    .C(_01437_),
    .X(_01439_));
 sky130_fd_sc_hd__and4_1 _10645_ (.A(net541),
    .B(net555),
    .C(net768),
    .D(net781),
    .X(_01440_));
 sky130_fd_sc_hd__a22oi_2 _10646_ (.A1(net555),
    .A2(net768),
    .B1(net781),
    .B2(net541),
    .Y(_01441_));
 sky130_fd_sc_hd__and4bb_1 _10647_ (.A_N(_01440_),
    .B_N(_01441_),
    .C(net572),
    .D(net757),
    .X(_01442_));
 sky130_fd_sc_hd__or2_2 _10648_ (.A(_01440_),
    .B(_01442_),
    .X(_01443_));
 sky130_fd_sc_hd__xnor2_4 _10649_ (.A(_01436_),
    .B(_01438_),
    .Y(_01444_));
 sky130_fd_sc_hd__nand2_2 _10650_ (.A(_01443_),
    .B(_01444_),
    .Y(_01445_));
 sky130_fd_sc_hd__a21oi_4 _10651_ (.A1(_01439_),
    .A2(_01445_),
    .B1(_01432_),
    .Y(_01446_));
 sky130_fd_sc_hd__a21o_1 _10652_ (.A1(_01439_),
    .A2(_01445_),
    .B1(_01432_),
    .X(_01447_));
 sky130_fd_sc_hd__nand3_2 _10653_ (.A(_01432_),
    .B(_01439_),
    .C(_01445_),
    .Y(_01448_));
 sky130_fd_sc_hd__o2bb2a_2 _10654_ (.A1_N(net599),
    .A2_N(net722),
    .B1(_01338_),
    .B2(_01339_),
    .X(_01449_));
 sky130_fd_sc_hd__nor2_4 _10655_ (.A(_01340_),
    .B(_01449_),
    .Y(_01450_));
 sky130_fd_sc_hd__and2_4 _10656_ (.A(net615),
    .B(net741),
    .X(_01451_));
 sky130_fd_sc_hd__and3_2 _10657_ (.A(net593),
    .B(net723),
    .C(_01451_),
    .X(_01452_));
 sky130_fd_sc_hd__a21oi_1 _10658_ (.A1(net587),
    .A2(net740),
    .B1(_01225_),
    .Y(_01453_));
 sky130_fd_sc_hd__and4bb_2 _10659_ (.A_N(_01452_),
    .B_N(_01453_),
    .C(net599),
    .D(net732),
    .X(_01454_));
 sky130_fd_sc_hd__nor2_4 _10660_ (.A(_01452_),
    .B(_01454_),
    .Y(_01455_));
 sky130_fd_sc_hd__xnor2_4 _10661_ (.A(_01450_),
    .B(_01455_),
    .Y(_01456_));
 sky130_fd_sc_hd__and3_4 _10662_ (.A(_01447_),
    .B(_01448_),
    .C(_01456_),
    .X(_01457_));
 sky130_fd_sc_hd__o211ai_4 _10663_ (.A1(_01446_),
    .A2(_01457_),
    .B1(_01430_),
    .C1(_01431_),
    .Y(_01458_));
 sky130_fd_sc_hd__a211o_1 _10664_ (.A1(_01430_),
    .A2(_01431_),
    .B1(_01446_),
    .C1(_01457_),
    .X(_01459_));
 sky130_fd_sc_hd__nand2_2 _10665_ (.A(_01458_),
    .B(_01459_),
    .Y(_01460_));
 sky130_fd_sc_hd__o211a_2 _10666_ (.A1(_01314_),
    .A2(_01383_),
    .B1(_01407_),
    .C1(_01427_),
    .X(_01461_));
 sky130_fd_sc_hd__nor3_4 _10667_ (.A(net120),
    .B(_01460_),
    .C(_01461_),
    .Y(_01462_));
 sky130_fd_sc_hd__o211ai_4 _10668_ (.A1(net120),
    .A2(_01462_),
    .B1(_01350_),
    .C1(_01382_),
    .Y(_01463_));
 sky130_fd_sc_hd__or3b_4 _10669_ (.A(_01354_),
    .B(_01455_),
    .C_N(_01450_),
    .X(_01464_));
 sky130_fd_sc_hd__nand2_4 _10670_ (.A(_01430_),
    .B(_01458_),
    .Y(_01465_));
 sky130_fd_sc_hd__nand2_1 _10671_ (.A(_01342_),
    .B(_01356_),
    .Y(_01466_));
 sky130_fd_sc_hd__and2_4 _10672_ (.A(_01357_),
    .B(_01466_),
    .X(_01467_));
 sky130_fd_sc_hd__xnor2_4 _10673_ (.A(_01465_),
    .B(_01467_),
    .Y(_01468_));
 sky130_fd_sc_hd__nor2_1 _10674_ (.A(_01464_),
    .B(_01468_),
    .Y(_01469_));
 sky130_fd_sc_hd__xor2_4 _10675_ (.A(_01464_),
    .B(_01468_),
    .X(_01470_));
 sky130_fd_sc_hd__a211o_2 _10676_ (.A1(_01350_),
    .A2(_01382_),
    .B1(net120),
    .C1(_01462_),
    .X(_01471_));
 sky130_fd_sc_hd__nand3_4 _10677_ (.A(_01463_),
    .B(_01470_),
    .C(_01471_),
    .Y(_01472_));
 sky130_fd_sc_hd__nand2_4 _10678_ (.A(_01463_),
    .B(_01472_),
    .Y(_01473_));
 sky130_fd_sc_hd__and2_2 _10679_ (.A(_01381_),
    .B(_01473_),
    .X(_01474_));
 sky130_fd_sc_hd__a21oi_4 _10680_ (.A1(_01465_),
    .A2(_01467_),
    .B1(_01469_),
    .Y(_01475_));
 sky130_fd_sc_hd__xnor2_4 _10681_ (.A(_01381_),
    .B(_01473_),
    .Y(_01476_));
 sky130_fd_sc_hd__nor2_2 _10682_ (.A(_01475_),
    .B(_01476_),
    .Y(_01477_));
 sky130_fd_sc_hd__o211ai_4 _10683_ (.A1(_01474_),
    .A2(_01477_),
    .B1(_01370_),
    .C1(_01380_),
    .Y(_01478_));
 sky130_fd_sc_hd__a211o_2 _10684_ (.A1(_01370_),
    .A2(_01380_),
    .B1(_01474_),
    .C1(_01477_),
    .X(_01479_));
 sky130_fd_sc_hd__nand3_4 _10685_ (.A(_01241_),
    .B(_01478_),
    .C(_01479_),
    .Y(_01480_));
 sky130_fd_sc_hd__o211a_2 _10686_ (.A1(_01373_),
    .A2(_01379_),
    .B1(_01478_),
    .C1(_01480_),
    .X(_01481_));
 sky130_fd_sc_hd__a21o_1 _10687_ (.A1(_01478_),
    .A2(_01479_),
    .B1(_01241_),
    .X(_01482_));
 sky130_fd_sc_hd__nand2_4 _10688_ (.A(_01480_),
    .B(_01482_),
    .Y(_01483_));
 sky130_fd_sc_hd__and2_1 _10689_ (.A(_01475_),
    .B(_01476_),
    .X(_01484_));
 sky130_fd_sc_hd__xor2_4 _10690_ (.A(_01475_),
    .B(_01476_),
    .X(_01485_));
 sky130_fd_sc_hd__a21o_1 _10691_ (.A1(_01463_),
    .A2(_01471_),
    .B1(_01470_),
    .X(_01486_));
 sky130_fd_sc_hd__o21a_2 _10692_ (.A1(net120),
    .A2(_01461_),
    .B1(_01460_),
    .X(_01487_));
 sky130_fd_sc_hd__a22oi_4 _10693_ (.A1(_01423_),
    .A2(_01424_),
    .B1(_01425_),
    .B2(_01407_),
    .Y(_01488_));
 sky130_fd_sc_hd__and4_1 _10694_ (.A(net431),
    .B(net440),
    .C(net903),
    .D(net918),
    .X(_01489_));
 sky130_fd_sc_hd__nand2_2 _10695_ (.A(net447),
    .B(net895),
    .Y(_01490_));
 sky130_fd_sc_hd__a22o_1 _10696_ (.A1(net440),
    .A2(net903),
    .B1(net918),
    .B2(net431),
    .X(_01491_));
 sky130_fd_sc_hd__and2b_2 _10697_ (.A_N(_01489_),
    .B(_01491_),
    .X(_01492_));
 sky130_fd_sc_hd__a31o_4 _10698_ (.A1(net447),
    .A2(net895),
    .A3(_01491_),
    .B1(_01489_),
    .X(_01493_));
 sky130_fd_sc_hd__xnor2_4 _10699_ (.A(_01400_),
    .B(_01402_),
    .Y(_01494_));
 sky130_fd_sc_hd__nand2_1 _10700_ (.A(_01493_),
    .B(_01494_),
    .Y(_01495_));
 sky130_fd_sc_hd__xor2_4 _10701_ (.A(_01493_),
    .B(_01494_),
    .X(_01496_));
 sky130_fd_sc_hd__and4_1 _10702_ (.A(net456),
    .B(net466),
    .C(net873),
    .D(net883),
    .X(_01497_));
 sky130_fd_sc_hd__nand2_4 _10703_ (.A(net475),
    .B(net864),
    .Y(_01498_));
 sky130_fd_sc_hd__a22oi_4 _10704_ (.A1(net466),
    .A2(net873),
    .B1(net883),
    .B2(net456),
    .Y(_01499_));
 sky130_fd_sc_hd__nor2_2 _10705_ (.A(_01497_),
    .B(_01499_),
    .Y(_01500_));
 sky130_fd_sc_hd__o21ba_2 _10706_ (.A1(_01498_),
    .A2(_01499_),
    .B1_N(_01497_),
    .X(_01501_));
 sky130_fd_sc_hd__nand2b_2 _10707_ (.A_N(_01501_),
    .B(_01496_),
    .Y(_01502_));
 sky130_fd_sc_hd__xnor2_4 _10708_ (.A(_01496_),
    .B(_01501_),
    .Y(_01503_));
 sky130_fd_sc_hd__xor2_4 _10709_ (.A(_01030_),
    .B(_01390_),
    .X(_01504_));
 sky130_fd_sc_hd__nand2_4 _10710_ (.A(_01503_),
    .B(_01504_),
    .Y(_01505_));
 sky130_fd_sc_hd__xnor2_4 _10711_ (.A(_01394_),
    .B(_01405_),
    .Y(_01506_));
 sky130_fd_sc_hd__or2_2 _10712_ (.A(_01505_),
    .B(_01506_),
    .X(_01507_));
 sky130_fd_sc_hd__xnor2_2 _10713_ (.A(_01419_),
    .B(_01421_),
    .Y(_01508_));
 sky130_fd_sc_hd__a21o_4 _10714_ (.A1(_01495_),
    .A2(_01502_),
    .B1(_01508_),
    .X(_01509_));
 sky130_fd_sc_hd__nand3_2 _10715_ (.A(_01495_),
    .B(_01502_),
    .C(_01508_),
    .Y(_01510_));
 sky130_fd_sc_hd__xnor2_4 _10716_ (.A(_01414_),
    .B(_01416_),
    .Y(_01511_));
 sky130_fd_sc_hd__and4_2 _10717_ (.A(net487),
    .B(net497),
    .C(net844),
    .D(net853),
    .X(_01512_));
 sky130_fd_sc_hd__a22oi_2 _10718_ (.A1(net497),
    .A2(net844),
    .B1(net853),
    .B2(net487),
    .Y(_01513_));
 sky130_fd_sc_hd__and4bb_4 _10719_ (.A_N(_01512_),
    .B_N(_01513_),
    .C(net504),
    .D(net834),
    .X(_01514_));
 sky130_fd_sc_hd__nor2_4 _10720_ (.A(_01512_),
    .B(_01514_),
    .Y(_01515_));
 sky130_fd_sc_hd__and2b_2 _10721_ (.A_N(_01515_),
    .B(_01511_),
    .X(_01516_));
 sky130_fd_sc_hd__xnor2_4 _10722_ (.A(_01511_),
    .B(_01515_),
    .Y(_01517_));
 sky130_fd_sc_hd__o2bb2a_1 _10723_ (.A1_N(net529),
    .A2_N(net791),
    .B1(_01433_),
    .B2(_01434_),
    .X(_01518_));
 sky130_fd_sc_hd__nor2_4 _10724_ (.A(_01435_),
    .B(_01518_),
    .Y(_01519_));
 sky130_fd_sc_hd__and2_2 _10725_ (.A(_01517_),
    .B(_01519_),
    .X(_01520_));
 sky130_fd_sc_hd__a211o_1 _10726_ (.A1(_01509_),
    .A2(_01510_),
    .B1(_01516_),
    .C1(_01520_),
    .X(_01521_));
 sky130_fd_sc_hd__o211ai_4 _10727_ (.A1(_01516_),
    .A2(_01520_),
    .B1(_01509_),
    .C1(_01510_),
    .Y(_01522_));
 sky130_fd_sc_hd__nand2_4 _10728_ (.A(_01521_),
    .B(_01522_),
    .Y(_01523_));
 sky130_fd_sc_hd__xor2_4 _10729_ (.A(_01505_),
    .B(_01506_),
    .X(_01524_));
 sky130_fd_sc_hd__nand2b_2 _10730_ (.A_N(_01523_),
    .B(_01524_),
    .Y(_01525_));
 sky130_fd_sc_hd__a211o_4 _10731_ (.A1(_01507_),
    .A2(_01525_),
    .B1(_01426_),
    .C1(_01488_),
    .X(_01526_));
 sky130_fd_sc_hd__a21oi_4 _10732_ (.A1(_01447_),
    .A2(_01448_),
    .B1(_01456_),
    .Y(_01527_));
 sky130_fd_sc_hd__a211oi_4 _10733_ (.A1(_01509_),
    .A2(_01522_),
    .B1(_01527_),
    .C1(_01457_),
    .Y(_01528_));
 sky130_fd_sc_hd__o211a_2 _10734_ (.A1(_01457_),
    .A2(_01527_),
    .B1(_01522_),
    .C1(_01509_),
    .X(_01529_));
 sky130_fd_sc_hd__xnor2_2 _10735_ (.A(_01443_),
    .B(_01444_),
    .Y(_01530_));
 sky130_fd_sc_hd__and4_2 _10736_ (.A(net513),
    .B(net520),
    .C(net814),
    .D(net825),
    .X(_01531_));
 sky130_fd_sc_hd__a22oi_2 _10737_ (.A1(net520),
    .A2(net814),
    .B1(net825),
    .B2(net513),
    .Y(_01532_));
 sky130_fd_sc_hd__and4bb_4 _10738_ (.A_N(_01531_),
    .B_N(_01532_),
    .C(net529),
    .D(net804),
    .X(_01533_));
 sky130_fd_sc_hd__nor2_4 _10739_ (.A(_01531_),
    .B(_01533_),
    .Y(_01534_));
 sky130_fd_sc_hd__o2bb2a_1 _10740_ (.A1_N(net572),
    .A2_N(net757),
    .B1(_01440_),
    .B2(_01441_),
    .X(_01535_));
 sky130_fd_sc_hd__nor2_2 _10741_ (.A(_01442_),
    .B(_01535_),
    .Y(_01536_));
 sky130_fd_sc_hd__or3_2 _10742_ (.A(_01442_),
    .B(_01534_),
    .C(_01535_),
    .X(_01537_));
 sky130_fd_sc_hd__and4_1 _10743_ (.A(net541),
    .B(net555),
    .C(net782),
    .D(net791),
    .X(_01538_));
 sky130_fd_sc_hd__a22oi_2 _10744_ (.A1(net555),
    .A2(net782),
    .B1(net791),
    .B2(net541),
    .Y(_01539_));
 sky130_fd_sc_hd__and4bb_1 _10745_ (.A_N(_01538_),
    .B_N(_01539_),
    .C(net572),
    .D(net768),
    .X(_01540_));
 sky130_fd_sc_hd__or2_2 _10746_ (.A(_01538_),
    .B(_01540_),
    .X(_01541_));
 sky130_fd_sc_hd__xnor2_4 _10747_ (.A(_01534_),
    .B(_01536_),
    .Y(_01542_));
 sky130_fd_sc_hd__nand2_1 _10748_ (.A(_01541_),
    .B(_01542_),
    .Y(_01543_));
 sky130_fd_sc_hd__a21o_4 _10749_ (.A1(_01537_),
    .A2(_01543_),
    .B1(_01530_),
    .X(_01544_));
 sky130_fd_sc_hd__nand3_2 _10750_ (.A(_01530_),
    .B(_01537_),
    .C(_01543_),
    .Y(_01545_));
 sky130_fd_sc_hd__o2bb2a_1 _10751_ (.A1_N(net599),
    .A2_N(net732),
    .B1(_01452_),
    .B2(_01453_),
    .X(_01546_));
 sky130_fd_sc_hd__and2_4 _10752_ (.A(net615),
    .B(net750),
    .X(_01547_));
 sky130_fd_sc_hd__and3_1 _10753_ (.A(net587),
    .B(net731),
    .C(_01547_),
    .X(_01548_));
 sky130_fd_sc_hd__a21oi_1 _10754_ (.A1(net587),
    .A2(net749),
    .B1(_01337_),
    .Y(_01549_));
 sky130_fd_sc_hd__and4bb_1 _10755_ (.A_N(_01548_),
    .B_N(_01549_),
    .C(net599),
    .D(net741),
    .X(_01550_));
 sky130_fd_sc_hd__nor2_1 _10756_ (.A(_01548_),
    .B(_01550_),
    .Y(_01551_));
 sky130_fd_sc_hd__or3_2 _10757_ (.A(_01454_),
    .B(_01546_),
    .C(_01551_),
    .X(_01552_));
 sky130_fd_sc_hd__o21ai_1 _10758_ (.A1(_01454_),
    .A2(_01546_),
    .B1(_01551_),
    .Y(_01553_));
 sky130_fd_sc_hd__and2_2 _10759_ (.A(_01552_),
    .B(_01553_),
    .X(_01554_));
 sky130_fd_sc_hd__and3_2 _10760_ (.A(_01544_),
    .B(_01545_),
    .C(_01554_),
    .X(_01555_));
 sky130_fd_sc_hd__inv_2 _10761_ (.A(_01555_),
    .Y(_01556_));
 sky130_fd_sc_hd__a211oi_4 _10762_ (.A1(_01544_),
    .A2(_01556_),
    .B1(_01528_),
    .C1(_01529_),
    .Y(_01557_));
 sky130_fd_sc_hd__o211a_1 _10763_ (.A1(_01528_),
    .A2(_01529_),
    .B1(_01544_),
    .C1(_01556_),
    .X(_01558_));
 sky130_fd_sc_hd__or2_1 _10764_ (.A(_01557_),
    .B(_01558_),
    .X(_01559_));
 sky130_fd_sc_hd__o211ai_4 _10765_ (.A1(_01426_),
    .A2(_01488_),
    .B1(_01507_),
    .C1(_01525_),
    .Y(_01560_));
 sky130_fd_sc_hd__nand3b_4 _10766_ (.A_N(_01559_),
    .B(_01560_),
    .C(_01526_),
    .Y(_01561_));
 sky130_fd_sc_hd__a211oi_4 _10767_ (.A1(_01526_),
    .A2(_01561_),
    .B1(_01462_),
    .C1(_01487_),
    .Y(_01562_));
 sky130_fd_sc_hd__o31ai_1 _10768_ (.A1(_01340_),
    .A2(_01449_),
    .A3(_01455_),
    .B1(_01354_),
    .Y(_01563_));
 sky130_fd_sc_hd__and2_1 _10769_ (.A(_01464_),
    .B(_01563_),
    .X(_01564_));
 sky130_fd_sc_hd__o21ai_2 _10770_ (.A1(_01528_),
    .A2(_01557_),
    .B1(_01564_),
    .Y(_01565_));
 sky130_fd_sc_hd__or3_1 _10771_ (.A(_01528_),
    .B(_01557_),
    .C(_01564_),
    .X(_01566_));
 sky130_fd_sc_hd__nand2_1 _10772_ (.A(_01565_),
    .B(_01566_),
    .Y(_01567_));
 sky130_fd_sc_hd__o211a_1 _10773_ (.A1(_01462_),
    .A2(_01487_),
    .B1(_01526_),
    .C1(_01561_),
    .X(_01568_));
 sky130_fd_sc_hd__nor3_2 _10774_ (.A(_01562_),
    .B(_01567_),
    .C(_01568_),
    .Y(_01569_));
 sky130_fd_sc_hd__o211a_2 _10775_ (.A1(_01562_),
    .A2(_01569_),
    .B1(_01472_),
    .C1(_01486_),
    .X(_01570_));
 sky130_fd_sc_hd__a211oi_2 _10776_ (.A1(_01472_),
    .A2(_01486_),
    .B1(_01562_),
    .C1(_01569_),
    .Y(_01571_));
 sky130_fd_sc_hd__nor3_2 _10777_ (.A(_01565_),
    .B(_01570_),
    .C(_01571_),
    .Y(_01572_));
 sky130_fd_sc_hd__nor2_4 _10778_ (.A(_01570_),
    .B(_01572_),
    .Y(_01573_));
 sky130_fd_sc_hd__xnor2_4 _10779_ (.A(_01485_),
    .B(_01573_),
    .Y(_01574_));
 sky130_fd_sc_hd__nand2_1 _10780_ (.A(_01355_),
    .B(_01574_),
    .Y(_01575_));
 sky130_fd_sc_hd__o31a_4 _10781_ (.A1(_01477_),
    .A2(_01484_),
    .A3(_01573_),
    .B1(_01575_),
    .X(_01576_));
 sky130_fd_sc_hd__a211oi_2 _10782_ (.A1(_01478_),
    .A2(_01480_),
    .B1(_01373_),
    .C1(_01379_),
    .Y(_01577_));
 sky130_fd_sc_hd__o21ba_1 _10783_ (.A1(_01483_),
    .A2(_01576_),
    .B1_N(_01577_),
    .X(_01578_));
 sky130_fd_sc_hd__xnor2_4 _10784_ (.A(_01483_),
    .B(_01576_),
    .Y(_01579_));
 sky130_fd_sc_hd__and2_4 _10785_ (.A(net612),
    .B(net758),
    .X(_01580_));
 sky130_fd_sc_hd__and3_1 _10786_ (.A(net588),
    .B(net782),
    .C(_01580_),
    .X(_01581_));
 sky130_fd_sc_hd__a21oi_1 _10787_ (.A1(net588),
    .A2(net782),
    .B1(_01580_),
    .Y(_01582_));
 sky130_fd_sc_hd__and4bb_2 _10788_ (.A_N(_01581_),
    .B_N(_01582_),
    .C(net600),
    .D(net769),
    .X(_01583_));
 sky130_fd_sc_hd__o2bb2a_1 _10789_ (.A1_N(net600),
    .A2_N(net769),
    .B1(_01581_),
    .B2(_01582_),
    .X(_01584_));
 sky130_fd_sc_hd__nor2_2 _10790_ (.A(_01583_),
    .B(_01584_),
    .Y(_01585_));
 sky130_fd_sc_hd__and4_1 _10791_ (.A(net588),
    .B(net612),
    .C(net771),
    .D(net792),
    .X(_01586_));
 sky130_fd_sc_hd__nand2_2 _10792_ (.A(net600),
    .B(net782),
    .Y(_01587_));
 sky130_fd_sc_hd__a22oi_4 _10793_ (.A1(net612),
    .A2(net771),
    .B1(net792),
    .B2(net588),
    .Y(_01588_));
 sky130_fd_sc_hd__nor2_1 _10794_ (.A(_01586_),
    .B(_01588_),
    .Y(_01589_));
 sky130_fd_sc_hd__o21ba_4 _10795_ (.A1(_01587_),
    .A2(_01588_),
    .B1_N(_01586_),
    .X(_01590_));
 sky130_fd_sc_hd__or3_4 _10796_ (.A(_01583_),
    .B(_01584_),
    .C(_01590_),
    .X(_01591_));
 sky130_fd_sc_hd__nand2_4 _10797_ (.A(net530),
    .B(net833),
    .Y(_01592_));
 sky130_fd_sc_hd__and2_2 _10798_ (.A(net522),
    .B(net847),
    .X(_01593_));
 sky130_fd_sc_hd__nand2_2 _10799_ (.A(net523),
    .B(net847),
    .Y(_01594_));
 sky130_fd_sc_hd__and3_1 _10800_ (.A(net512),
    .B(net859),
    .C(_01593_),
    .X(_01595_));
 sky130_fd_sc_hd__a21oi_2 _10801_ (.A1(net512),
    .A2(net853),
    .B1(_01593_),
    .Y(_01596_));
 sky130_fd_sc_hd__nor2_2 _10802_ (.A(_01595_),
    .B(_01596_),
    .Y(_01597_));
 sky130_fd_sc_hd__xnor2_4 _10803_ (.A(_01592_),
    .B(_01597_),
    .Y(_01598_));
 sky130_fd_sc_hd__nand2_4 _10804_ (.A(net504),
    .B(net864),
    .Y(_01599_));
 sky130_fd_sc_hd__and4_1 _10805_ (.A(net486),
    .B(net496),
    .C(net873),
    .D(net884),
    .X(_01600_));
 sky130_fd_sc_hd__a22oi_4 _10806_ (.A1(net496),
    .A2(net874),
    .B1(net884),
    .B2(net486),
    .Y(_01601_));
 sky130_fd_sc_hd__nor2_2 _10807_ (.A(_01600_),
    .B(_01601_),
    .Y(_01602_));
 sky130_fd_sc_hd__xnor2_4 _10808_ (.A(_01599_),
    .B(_01602_),
    .Y(_01603_));
 sky130_fd_sc_hd__and4_1 _10809_ (.A(net486),
    .B(net496),
    .C(net884),
    .D(net895),
    .X(_01604_));
 sky130_fd_sc_hd__a22oi_2 _10810_ (.A1(net496),
    .A2(net883),
    .B1(net895),
    .B2(net486),
    .Y(_01605_));
 sky130_fd_sc_hd__and4bb_2 _10811_ (.A_N(_01604_),
    .B_N(_01605_),
    .C(net504),
    .D(net873),
    .X(_01606_));
 sky130_fd_sc_hd__nor2_2 _10812_ (.A(_01604_),
    .B(_01606_),
    .Y(_01607_));
 sky130_fd_sc_hd__nand2b_1 _10813_ (.A_N(_01607_),
    .B(_01603_),
    .Y(_01608_));
 sky130_fd_sc_hd__xnor2_2 _10814_ (.A(_01603_),
    .B(_01607_),
    .Y(_01609_));
 sky130_fd_sc_hd__nand2_1 _10815_ (.A(_01598_),
    .B(_01609_),
    .Y(_01610_));
 sky130_fd_sc_hd__xnor2_1 _10816_ (.A(_01598_),
    .B(_01609_),
    .Y(_01611_));
 sky130_fd_sc_hd__o2bb2a_1 _10817_ (.A1_N(net504),
    .A2_N(net873),
    .B1(_01604_),
    .B2(_01605_),
    .X(_01612_));
 sky130_fd_sc_hd__nor2_1 _10818_ (.A(_01606_),
    .B(_01612_),
    .Y(_01613_));
 sky130_fd_sc_hd__and4_1 _10819_ (.A(net488),
    .B(net498),
    .C(net896),
    .D(net908),
    .X(_01614_));
 sky130_fd_sc_hd__a22oi_2 _10820_ (.A1(net498),
    .A2(net895),
    .B1(net908),
    .B2(net488),
    .Y(_01615_));
 sky130_fd_sc_hd__and4bb_2 _10821_ (.A_N(_01614_),
    .B_N(_01615_),
    .C(net505),
    .D(net888),
    .X(_01616_));
 sky130_fd_sc_hd__nor2_2 _10822_ (.A(_01614_),
    .B(_01616_),
    .Y(_01617_));
 sky130_fd_sc_hd__or3_1 _10823_ (.A(_01606_),
    .B(_01612_),
    .C(_01617_),
    .X(_01618_));
 sky130_fd_sc_hd__nand2_4 _10824_ (.A(net530),
    .B(net846),
    .Y(_01619_));
 sky130_fd_sc_hd__and4_1 _10825_ (.A(net512),
    .B(net524),
    .C(net856),
    .D(net865),
    .X(_01620_));
 sky130_fd_sc_hd__a22oi_4 _10826_ (.A1(net521),
    .A2(net856),
    .B1(net866),
    .B2(net512),
    .Y(_01621_));
 sky130_fd_sc_hd__nor2_2 _10827_ (.A(_01620_),
    .B(_01621_),
    .Y(_01622_));
 sky130_fd_sc_hd__xnor2_4 _10828_ (.A(_01619_),
    .B(_01622_),
    .Y(_01623_));
 sky130_fd_sc_hd__xnor2_2 _10829_ (.A(_01613_),
    .B(_01617_),
    .Y(_01624_));
 sky130_fd_sc_hd__nand2_1 _10830_ (.A(_01623_),
    .B(_01624_),
    .Y(_01625_));
 sky130_fd_sc_hd__a21o_2 _10831_ (.A1(_01618_),
    .A2(_01625_),
    .B1(_01611_),
    .X(_01626_));
 sky130_fd_sc_hd__inv_2 _10832_ (.A(_01626_),
    .Y(_01627_));
 sky130_fd_sc_hd__and4_1 _10833_ (.A(net542),
    .B(net556),
    .C(net820),
    .D(net828),
    .X(_01628_));
 sky130_fd_sc_hd__a22oi_2 _10834_ (.A1(net556),
    .A2(net820),
    .B1(net828),
    .B2(net542),
    .Y(_01629_));
 sky130_fd_sc_hd__and4bb_2 _10835_ (.A_N(_01628_),
    .B_N(_01629_),
    .C(net573),
    .D(net804),
    .X(_01630_));
 sky130_fd_sc_hd__or2_4 _10836_ (.A(_01628_),
    .B(_01630_),
    .X(_01631_));
 sky130_fd_sc_hd__o21ba_2 _10837_ (.A1(_01592_),
    .A2(_01596_),
    .B1_N(_01595_),
    .X(_01632_));
 sky130_fd_sc_hd__nand2_2 _10838_ (.A(net573),
    .B(net792),
    .Y(_01633_));
 sky130_fd_sc_hd__and4_2 _10839_ (.A(net542),
    .B(net556),
    .C(net805),
    .D(net820),
    .X(_01634_));
 sky130_fd_sc_hd__a22oi_4 _10840_ (.A1(net556),
    .A2(net805),
    .B1(net820),
    .B2(net542),
    .Y(_01635_));
 sky130_fd_sc_hd__nor2_4 _10841_ (.A(_01634_),
    .B(_01635_),
    .Y(_01636_));
 sky130_fd_sc_hd__xnor2_4 _10842_ (.A(_01633_),
    .B(_01636_),
    .Y(_01637_));
 sky130_fd_sc_hd__nand2b_2 _10843_ (.A_N(_01632_),
    .B(_01637_),
    .Y(_01638_));
 sky130_fd_sc_hd__xnor2_4 _10844_ (.A(_01632_),
    .B(_01637_),
    .Y(_01639_));
 sky130_fd_sc_hd__nand2_2 _10845_ (.A(_01631_),
    .B(_01639_),
    .Y(_01640_));
 sky130_fd_sc_hd__xnor2_4 _10846_ (.A(_01631_),
    .B(_01639_),
    .Y(_01641_));
 sky130_fd_sc_hd__o21ba_4 _10847_ (.A1(_01619_),
    .A2(_01621_),
    .B1_N(_01620_),
    .X(_01642_));
 sky130_fd_sc_hd__o22a_1 _10848_ (.A1(net303),
    .A2(_03269_),
    .B1(_01628_),
    .B2(_01629_),
    .X(_01643_));
 sky130_fd_sc_hd__nor2_2 _10849_ (.A(_01630_),
    .B(_01643_),
    .Y(_01644_));
 sky130_fd_sc_hd__or3_4 _10850_ (.A(_01630_),
    .B(_01642_),
    .C(_01643_),
    .X(_01645_));
 sky130_fd_sc_hd__and4_1 _10851_ (.A(net542),
    .B(net556),
    .C(net828),
    .D(net835),
    .X(_01646_));
 sky130_fd_sc_hd__a22oi_2 _10852_ (.A1(net561),
    .A2(net828),
    .B1(net835),
    .B2(net542),
    .Y(_01647_));
 sky130_fd_sc_hd__and4bb_2 _10853_ (.A_N(_01646_),
    .B_N(_01647_),
    .C(net573),
    .D(net817),
    .X(_01648_));
 sky130_fd_sc_hd__or2_4 _10854_ (.A(_01646_),
    .B(_01648_),
    .X(_01649_));
 sky130_fd_sc_hd__xnor2_4 _10855_ (.A(_01642_),
    .B(_01644_),
    .Y(_01650_));
 sky130_fd_sc_hd__nand2_2 _10856_ (.A(_01649_),
    .B(_01650_),
    .Y(_01651_));
 sky130_fd_sc_hd__a21oi_4 _10857_ (.A1(_01645_),
    .A2(_01651_),
    .B1(_01641_),
    .Y(_01652_));
 sky130_fd_sc_hd__a21o_1 _10858_ (.A1(_01645_),
    .A2(_01651_),
    .B1(_01641_),
    .X(_01653_));
 sky130_fd_sc_hd__nand3_2 _10859_ (.A(_01641_),
    .B(_01645_),
    .C(_01651_),
    .Y(_01654_));
 sky130_fd_sc_hd__xnor2_4 _10860_ (.A(_01585_),
    .B(_01590_),
    .Y(_01655_));
 sky130_fd_sc_hd__and3_4 _10861_ (.A(_01653_),
    .B(_01654_),
    .C(_01655_),
    .X(_01656_));
 sky130_fd_sc_hd__a21oi_4 _10862_ (.A1(_01653_),
    .A2(_01654_),
    .B1(_01655_),
    .Y(_01657_));
 sky130_fd_sc_hd__or3_4 _10863_ (.A(_01626_),
    .B(_01656_),
    .C(_01657_),
    .X(_01658_));
 sky130_fd_sc_hd__o21ai_4 _10864_ (.A1(_01656_),
    .A2(_01657_),
    .B1(_01626_),
    .Y(_01659_));
 sky130_fd_sc_hd__xnor2_4 _10865_ (.A(_01649_),
    .B(_01650_),
    .Y(_01660_));
 sky130_fd_sc_hd__and4_4 _10866_ (.A(net512),
    .B(net522),
    .C(net865),
    .D(net876),
    .X(_01661_));
 sky130_fd_sc_hd__and2_2 _10867_ (.A(net532),
    .B(net857),
    .X(_01662_));
 sky130_fd_sc_hd__nand2_4 _10868_ (.A(net532),
    .B(net857),
    .Y(_01663_));
 sky130_fd_sc_hd__a22oi_4 _10869_ (.A1(net522),
    .A2(net865),
    .B1(net876),
    .B2(net512),
    .Y(_01664_));
 sky130_fd_sc_hd__nor2_4 _10870_ (.A(_01661_),
    .B(_01664_),
    .Y(_01665_));
 sky130_fd_sc_hd__a21oi_4 _10871_ (.A1(_01662_),
    .A2(_01665_),
    .B1(_01661_),
    .Y(_01666_));
 sky130_fd_sc_hd__o2bb2a_1 _10872_ (.A1_N(net573),
    .A2_N(net817),
    .B1(_01646_),
    .B2(_01647_),
    .X(_01667_));
 sky130_fd_sc_hd__nor2_2 _10873_ (.A(_01648_),
    .B(_01667_),
    .Y(_01668_));
 sky130_fd_sc_hd__or3_4 _10874_ (.A(_01648_),
    .B(_01666_),
    .C(_01667_),
    .X(_01669_));
 sky130_fd_sc_hd__and4_1 _10875_ (.A(net542),
    .B(net556),
    .C(net835),
    .D(net846),
    .X(_01670_));
 sky130_fd_sc_hd__a22oi_2 _10876_ (.A1(net556),
    .A2(net835),
    .B1(net846),
    .B2(net542),
    .Y(_01671_));
 sky130_fd_sc_hd__and4bb_2 _10877_ (.A_N(_01670_),
    .B_N(_01671_),
    .C(net573),
    .D(net825),
    .X(_01672_));
 sky130_fd_sc_hd__or2_4 _10878_ (.A(_01670_),
    .B(_01672_),
    .X(_01673_));
 sky130_fd_sc_hd__xnor2_4 _10879_ (.A(_01666_),
    .B(_01668_),
    .Y(_01674_));
 sky130_fd_sc_hd__nand2_2 _10880_ (.A(_01673_),
    .B(_01674_),
    .Y(_01675_));
 sky130_fd_sc_hd__a21oi_4 _10881_ (.A1(_01669_),
    .A2(_01675_),
    .B1(_01660_),
    .Y(_01676_));
 sky130_fd_sc_hd__a21o_1 _10882_ (.A1(_01669_),
    .A2(_01675_),
    .B1(_01660_),
    .X(_01677_));
 sky130_fd_sc_hd__nand3_2 _10883_ (.A(_01660_),
    .B(_01669_),
    .C(_01675_),
    .Y(_01678_));
 sky130_fd_sc_hd__xnor2_2 _10884_ (.A(_01587_),
    .B(_01589_),
    .Y(_01679_));
 sky130_fd_sc_hd__and4_4 _10885_ (.A(net588),
    .B(net612),
    .C(net782),
    .D(net805),
    .X(_01680_));
 sky130_fd_sc_hd__nand2_2 _10886_ (.A(net602),
    .B(net792),
    .Y(_01681_));
 sky130_fd_sc_hd__o2bb2a_2 _10887_ (.A1_N(net612),
    .A2_N(net782),
    .B1(_03269_),
    .B2(_03225_),
    .X(_01682_));
 sky130_fd_sc_hd__nor2_4 _10888_ (.A(_01680_),
    .B(_01682_),
    .Y(_01683_));
 sky130_fd_sc_hd__and3_2 _10889_ (.A(net600),
    .B(net792),
    .C(_01683_),
    .X(_01684_));
 sky130_fd_sc_hd__o21ai_4 _10890_ (.A1(_01680_),
    .A2(_01684_),
    .B1(_01679_),
    .Y(_01685_));
 sky130_fd_sc_hd__or3_1 _10891_ (.A(_01679_),
    .B(_01680_),
    .C(_01684_),
    .X(_01686_));
 sky130_fd_sc_hd__and2_2 _10892_ (.A(_01685_),
    .B(_01686_),
    .X(_01687_));
 sky130_fd_sc_hd__and3_4 _10893_ (.A(_01677_),
    .B(_01678_),
    .C(_01687_),
    .X(_01688_));
 sky130_fd_sc_hd__o211ai_4 _10894_ (.A1(_01676_),
    .A2(_01688_),
    .B1(_01658_),
    .C1(_01659_),
    .Y(_01689_));
 sky130_fd_sc_hd__and2_2 _10895_ (.A(_01658_),
    .B(_01689_),
    .X(_01690_));
 sky130_fd_sc_hd__or2_4 _10896_ (.A(_01591_),
    .B(_01690_),
    .X(_01691_));
 sky130_fd_sc_hd__and3_1 _10897_ (.A(net588),
    .B(net769),
    .C(_01547_),
    .X(_01692_));
 sky130_fd_sc_hd__a21oi_1 _10898_ (.A1(net588),
    .A2(net769),
    .B1(_01547_),
    .Y(_01693_));
 sky130_fd_sc_hd__and4bb_1 _10899_ (.A_N(_01692_),
    .B_N(_01693_),
    .C(net605),
    .D(net758),
    .X(_01694_));
 sky130_fd_sc_hd__o2bb2a_1 _10900_ (.A1_N(net605),
    .A2_N(net758),
    .B1(_01692_),
    .B2(_01693_),
    .X(_01695_));
 sky130_fd_sc_hd__nor2_1 _10901_ (.A(_01581_),
    .B(_01583_),
    .Y(_01696_));
 sky130_fd_sc_hd__or3_4 _10902_ (.A(_01694_),
    .B(_01695_),
    .C(_01696_),
    .X(_01697_));
 sky130_fd_sc_hd__nand2_1 _10903_ (.A(net476),
    .B(net916),
    .Y(_01698_));
 sky130_fd_sc_hd__and4_1 _10904_ (.A(net466),
    .B(net475),
    .C(net903),
    .D(net913),
    .X(_01699_));
 sky130_fd_sc_hd__and4_1 _10905_ (.A(net456),
    .B(net468),
    .C(net903),
    .D(net913),
    .X(_01700_));
 sky130_fd_sc_hd__a22oi_2 _10906_ (.A1(net467),
    .A2(net904),
    .B1(net913),
    .B2(net456),
    .Y(_01701_));
 sky130_fd_sc_hd__nor2_1 _10907_ (.A(_01700_),
    .B(_01701_),
    .Y(_01702_));
 sky130_fd_sc_hd__nand2_2 _10908_ (.A(net475),
    .B(net896),
    .Y(_01703_));
 sky130_fd_sc_hd__xnor2_2 _10909_ (.A(_01702_),
    .B(_01703_),
    .Y(_01704_));
 sky130_fd_sc_hd__nand2_2 _10910_ (.A(_01699_),
    .B(_01704_),
    .Y(_01705_));
 sky130_fd_sc_hd__nand2_4 _10911_ (.A(net504),
    .B(net859),
    .Y(_01706_));
 sky130_fd_sc_hd__and4_1 _10912_ (.A(net486),
    .B(net497),
    .C(net864),
    .D(net874),
    .X(_01707_));
 sky130_fd_sc_hd__a22oi_4 _10913_ (.A1(net496),
    .A2(net864),
    .B1(net874),
    .B2(net487),
    .Y(_01708_));
 sky130_fd_sc_hd__nor2_2 _10914_ (.A(_01707_),
    .B(_01708_),
    .Y(_01709_));
 sky130_fd_sc_hd__xnor2_4 _10915_ (.A(_01706_),
    .B(_01709_),
    .Y(_01710_));
 sky130_fd_sc_hd__o21ba_1 _10916_ (.A1(_01599_),
    .A2(_01601_),
    .B1_N(_01600_),
    .X(_01711_));
 sky130_fd_sc_hd__and2b_1 _10917_ (.A_N(_01711_),
    .B(_01710_),
    .X(_01712_));
 sky130_fd_sc_hd__xnor2_2 _10918_ (.A(_01710_),
    .B(_01711_),
    .Y(_01713_));
 sky130_fd_sc_hd__nand2_2 _10919_ (.A(net531),
    .B(net827),
    .Y(_01714_));
 sky130_fd_sc_hd__and2_4 _10920_ (.A(net512),
    .B(net836),
    .X(_01715_));
 sky130_fd_sc_hd__nand2_1 _10921_ (.A(net514),
    .B(net836),
    .Y(_01716_));
 sky130_fd_sc_hd__a22o_1 _10922_ (.A1(net522),
    .A2(net836),
    .B1(net847),
    .B2(net512),
    .X(_01717_));
 sky130_fd_sc_hd__o21a_2 _10923_ (.A1(_01594_),
    .A2(_01716_),
    .B1(_01717_),
    .X(_01718_));
 sky130_fd_sc_hd__xnor2_4 _10924_ (.A(_01714_),
    .B(_01718_),
    .Y(_01719_));
 sky130_fd_sc_hd__and2_1 _10925_ (.A(_01713_),
    .B(_01719_),
    .X(_01720_));
 sky130_fd_sc_hd__xnor2_2 _10926_ (.A(_01713_),
    .B(_01719_),
    .Y(_01721_));
 sky130_fd_sc_hd__or2_2 _10927_ (.A(_01705_),
    .B(_01721_),
    .X(_01722_));
 sky130_fd_sc_hd__xnor2_2 _10928_ (.A(_01705_),
    .B(_01721_),
    .Y(_01723_));
 sky130_fd_sc_hd__a21o_4 _10929_ (.A1(_01608_),
    .A2(_01610_),
    .B1(_01723_),
    .X(_01724_));
 sky130_fd_sc_hd__a31o_4 _10930_ (.A1(net573),
    .A2(net792),
    .A3(_01636_),
    .B1(_01634_),
    .X(_01725_));
 sky130_fd_sc_hd__a32o_4 _10931_ (.A1(net530),
    .A2(net827),
    .A3(_01717_),
    .B1(_01715_),
    .B2(_01593_),
    .X(_01726_));
 sky130_fd_sc_hd__nand2_2 _10932_ (.A(net572),
    .B(net781),
    .Y(_01727_));
 sky130_fd_sc_hd__and4_2 _10933_ (.A(net541),
    .B(net555),
    .C(net791),
    .D(net804),
    .X(_01728_));
 sky130_fd_sc_hd__a22oi_4 _10934_ (.A1(net555),
    .A2(net794),
    .B1(net805),
    .B2(net541),
    .Y(_01729_));
 sky130_fd_sc_hd__nor2_4 _10935_ (.A(_01728_),
    .B(_01729_),
    .Y(_01730_));
 sky130_fd_sc_hd__xnor2_4 _10936_ (.A(_01727_),
    .B(_01730_),
    .Y(_01731_));
 sky130_fd_sc_hd__nand2_2 _10937_ (.A(_01726_),
    .B(_01731_),
    .Y(_01732_));
 sky130_fd_sc_hd__xor2_4 _10938_ (.A(_01726_),
    .B(_01731_),
    .X(_01733_));
 sky130_fd_sc_hd__nand2_2 _10939_ (.A(_01725_),
    .B(_01733_),
    .Y(_01734_));
 sky130_fd_sc_hd__xnor2_4 _10940_ (.A(_01725_),
    .B(_01733_),
    .Y(_01735_));
 sky130_fd_sc_hd__a21oi_4 _10941_ (.A1(_01638_),
    .A2(_01640_),
    .B1(_01735_),
    .Y(_01736_));
 sky130_fd_sc_hd__a21o_1 _10942_ (.A1(_01638_),
    .A2(_01640_),
    .B1(_01735_),
    .X(_01737_));
 sky130_fd_sc_hd__nand3_2 _10943_ (.A(_01638_),
    .B(_01640_),
    .C(_01735_),
    .Y(_01738_));
 sky130_fd_sc_hd__o21ai_1 _10944_ (.A1(_01694_),
    .A2(_01695_),
    .B1(_01696_),
    .Y(_01739_));
 sky130_fd_sc_hd__and2_2 _10945_ (.A(_01697_),
    .B(_01739_),
    .X(_01740_));
 sky130_fd_sc_hd__and3_4 _10946_ (.A(_01737_),
    .B(_01738_),
    .C(_01740_),
    .X(_01741_));
 sky130_fd_sc_hd__a21oi_4 _10947_ (.A1(_01737_),
    .A2(_01738_),
    .B1(_01740_),
    .Y(_01742_));
 sky130_fd_sc_hd__a211o_2 _10948_ (.A1(_01722_),
    .A2(_01724_),
    .B1(_01741_),
    .C1(_01742_),
    .X(_01743_));
 sky130_fd_sc_hd__o211ai_4 _10949_ (.A1(_01741_),
    .A2(_01742_),
    .B1(_01722_),
    .C1(_01724_),
    .Y(_01744_));
 sky130_fd_sc_hd__o211ai_4 _10950_ (.A1(_01652_),
    .A2(_01656_),
    .B1(_01743_),
    .C1(_01744_),
    .Y(_01745_));
 sky130_fd_sc_hd__and2_2 _10951_ (.A(_01743_),
    .B(_01745_),
    .X(_01746_));
 sky130_fd_sc_hd__or2_4 _10952_ (.A(_01697_),
    .B(_01746_),
    .X(_01747_));
 sky130_fd_sc_hd__xnor2_4 _10953_ (.A(_01697_),
    .B(_01746_),
    .Y(_01748_));
 sky130_fd_sc_hd__and4_1 _10954_ (.A(net457),
    .B(net468),
    .C(net895),
    .D(net903),
    .X(_01749_));
 sky130_fd_sc_hd__inv_2 _10955_ (.A(_01749_),
    .Y(_01750_));
 sky130_fd_sc_hd__a22o_2 _10956_ (.A1(net468),
    .A2(net895),
    .B1(net904),
    .B2(net458),
    .X(_01751_));
 sky130_fd_sc_hd__and4b_2 _10957_ (.A_N(_01749_),
    .B(_01751_),
    .C(net476),
    .D(net884),
    .X(_01752_));
 sky130_fd_sc_hd__a22oi_4 _10958_ (.A1(net476),
    .A2(net884),
    .B1(_01750_),
    .B2(_01751_),
    .Y(_01753_));
 sky130_fd_sc_hd__nor2_2 _10959_ (.A(_01752_),
    .B(_01753_),
    .Y(_01754_));
 sky130_fd_sc_hd__o21ba_2 _10960_ (.A1(_01701_),
    .A2(_01703_),
    .B1_N(_01700_),
    .X(_01755_));
 sky130_fd_sc_hd__or3_4 _10961_ (.A(_01752_),
    .B(_01753_),
    .C(_01755_),
    .X(_01756_));
 sky130_fd_sc_hd__nand2_4 _10962_ (.A(net504),
    .B(net844),
    .Y(_01757_));
 sky130_fd_sc_hd__and4_1 _10963_ (.A(net487),
    .B(net497),
    .C(net853),
    .D(net864),
    .X(_01758_));
 sky130_fd_sc_hd__a22oi_4 _10964_ (.A1(net497),
    .A2(net853),
    .B1(net864),
    .B2(net487),
    .Y(_01759_));
 sky130_fd_sc_hd__nor2_2 _10965_ (.A(_01758_),
    .B(_01759_),
    .Y(_01760_));
 sky130_fd_sc_hd__xnor2_4 _10966_ (.A(_01757_),
    .B(_01760_),
    .Y(_01761_));
 sky130_fd_sc_hd__o21ba_2 _10967_ (.A1(_01706_),
    .A2(_01708_),
    .B1_N(_01707_),
    .X(_01762_));
 sky130_fd_sc_hd__and2b_2 _10968_ (.A_N(_01762_),
    .B(_01761_),
    .X(_01763_));
 sky130_fd_sc_hd__xnor2_4 _10969_ (.A(_01761_),
    .B(_01762_),
    .Y(_01764_));
 sky130_fd_sc_hd__nand2_4 _10970_ (.A(net529),
    .B(net814),
    .Y(_01765_));
 sky130_fd_sc_hd__and3_1 _10971_ (.A(net520),
    .B(net826),
    .C(_01715_),
    .X(_01766_));
 sky130_fd_sc_hd__a21oi_2 _10972_ (.A1(net520),
    .A2(net825),
    .B1(_01715_),
    .Y(_01767_));
 sky130_fd_sc_hd__nor2_2 _10973_ (.A(_01766_),
    .B(_01767_),
    .Y(_01768_));
 sky130_fd_sc_hd__xnor2_4 _10974_ (.A(_01765_),
    .B(_01768_),
    .Y(_01769_));
 sky130_fd_sc_hd__and2_1 _10975_ (.A(_01764_),
    .B(_01769_),
    .X(_01770_));
 sky130_fd_sc_hd__xnor2_4 _10976_ (.A(_01764_),
    .B(_01769_),
    .Y(_01771_));
 sky130_fd_sc_hd__or2_2 _10977_ (.A(_01756_),
    .B(_01771_),
    .X(_01772_));
 sky130_fd_sc_hd__xor2_4 _10978_ (.A(_01756_),
    .B(_01771_),
    .X(_01773_));
 sky130_fd_sc_hd__o21ai_4 _10979_ (.A1(_01712_),
    .A2(_01720_),
    .B1(_01773_),
    .Y(_01774_));
 sky130_fd_sc_hd__a31o_4 _10980_ (.A1(net572),
    .A2(net781),
    .A3(_01730_),
    .B1(_01728_),
    .X(_01775_));
 sky130_fd_sc_hd__o21ba_4 _10981_ (.A1(_01765_),
    .A2(_01767_),
    .B1_N(_01766_),
    .X(_01776_));
 sky130_fd_sc_hd__o2bb2a_1 _10982_ (.A1_N(net572),
    .A2_N(net768),
    .B1(_01538_),
    .B2(_01539_),
    .X(_01777_));
 sky130_fd_sc_hd__nor2_2 _10983_ (.A(_01540_),
    .B(_01777_),
    .Y(_01778_));
 sky130_fd_sc_hd__or3_2 _10984_ (.A(_01540_),
    .B(_01776_),
    .C(_01777_),
    .X(_01779_));
 sky130_fd_sc_hd__xnor2_4 _10985_ (.A(_01776_),
    .B(_01778_),
    .Y(_01780_));
 sky130_fd_sc_hd__nand2_2 _10986_ (.A(_01775_),
    .B(_01780_),
    .Y(_01781_));
 sky130_fd_sc_hd__xnor2_4 _10987_ (.A(_01775_),
    .B(_01780_),
    .Y(_01782_));
 sky130_fd_sc_hd__a21oi_4 _10988_ (.A1(_01732_),
    .A2(_01734_),
    .B1(_01782_),
    .Y(_01783_));
 sky130_fd_sc_hd__a21o_1 _10989_ (.A1(_01732_),
    .A2(_01734_),
    .B1(_01782_),
    .X(_01784_));
 sky130_fd_sc_hd__nand3_2 _10990_ (.A(_01732_),
    .B(_01734_),
    .C(_01782_),
    .Y(_01785_));
 sky130_fd_sc_hd__and3_1 _10991_ (.A(net588),
    .B(net740),
    .C(_01580_),
    .X(_01786_));
 sky130_fd_sc_hd__a21oi_1 _10992_ (.A1(net588),
    .A2(net758),
    .B1(_01451_),
    .Y(_01787_));
 sky130_fd_sc_hd__and4bb_1 _10993_ (.A_N(_01786_),
    .B_N(_01787_),
    .C(net605),
    .D(net749),
    .X(_01788_));
 sky130_fd_sc_hd__o2bb2a_1 _10994_ (.A1_N(net600),
    .A2_N(net749),
    .B1(_01786_),
    .B2(_01787_),
    .X(_01789_));
 sky130_fd_sc_hd__nor2_1 _10995_ (.A(_01692_),
    .B(_01694_),
    .Y(_01790_));
 sky130_fd_sc_hd__or3_4 _10996_ (.A(_01788_),
    .B(_01789_),
    .C(_01790_),
    .X(_01791_));
 sky130_fd_sc_hd__o21ai_1 _10997_ (.A1(_01788_),
    .A2(_01789_),
    .B1(_01790_),
    .Y(_01792_));
 sky130_fd_sc_hd__and2_2 _10998_ (.A(_01791_),
    .B(_01792_),
    .X(_01793_));
 sky130_fd_sc_hd__and3_4 _10999_ (.A(_01784_),
    .B(_01785_),
    .C(_01793_),
    .X(_01794_));
 sky130_fd_sc_hd__a21oi_4 _11000_ (.A1(_01784_),
    .A2(_01785_),
    .B1(_01793_),
    .Y(_01795_));
 sky130_fd_sc_hd__a211o_2 _11001_ (.A1(_01772_),
    .A2(_01774_),
    .B1(_01794_),
    .C1(_01795_),
    .X(_01796_));
 sky130_fd_sc_hd__o211ai_4 _11002_ (.A1(_01794_),
    .A2(_01795_),
    .B1(_01772_),
    .C1(_01774_),
    .Y(_01797_));
 sky130_fd_sc_hd__o211ai_4 _11003_ (.A1(_01736_),
    .A2(_01741_),
    .B1(_01796_),
    .C1(_01797_),
    .Y(_01798_));
 sky130_fd_sc_hd__a211o_2 _11004_ (.A1(_01796_),
    .A2(_01797_),
    .B1(_01736_),
    .C1(_01741_),
    .X(_01799_));
 sky130_fd_sc_hd__nand2_2 _11005_ (.A(net476),
    .B(net873),
    .Y(_01800_));
 sky130_fd_sc_hd__and3_1 _11006_ (.A(net456),
    .B(net466),
    .C(net894),
    .X(_01801_));
 sky130_fd_sc_hd__a22o_1 _11007_ (.A1(net466),
    .A2(net883),
    .B1(net894),
    .B2(net456),
    .X(_01802_));
 sky130_fd_sc_hd__a21bo_2 _11008_ (.A1(net883),
    .A2(_01801_),
    .B1_N(_01802_),
    .X(_01803_));
 sky130_fd_sc_hd__xor2_4 _11009_ (.A(_01800_),
    .B(_01803_),
    .X(_01804_));
 sky130_fd_sc_hd__nor2_1 _11010_ (.A(_01749_),
    .B(_01752_),
    .Y(_01805_));
 sky130_fd_sc_hd__nand2b_4 _11011_ (.A_N(_01805_),
    .B(_01804_),
    .Y(_01806_));
 sky130_fd_sc_hd__o2bb2a_1 _11012_ (.A1_N(net504),
    .A2_N(net834),
    .B1(_01512_),
    .B2(_01513_),
    .X(_01807_));
 sky130_fd_sc_hd__nor2_4 _11013_ (.A(_01514_),
    .B(_01807_),
    .Y(_01808_));
 sky130_fd_sc_hd__o21ba_2 _11014_ (.A1(_01757_),
    .A2(_01759_),
    .B1_N(_01758_),
    .X(_01809_));
 sky130_fd_sc_hd__and2b_4 _11015_ (.A_N(_01809_),
    .B(_01808_),
    .X(_01810_));
 sky130_fd_sc_hd__xnor2_4 _11016_ (.A(_01808_),
    .B(_01809_),
    .Y(_01811_));
 sky130_fd_sc_hd__o2bb2a_1 _11017_ (.A1_N(net529),
    .A2_N(net804),
    .B1(_01531_),
    .B2(_01532_),
    .X(_01812_));
 sky130_fd_sc_hd__nor2_4 _11018_ (.A(_01533_),
    .B(_01812_),
    .Y(_01813_));
 sky130_fd_sc_hd__and2_2 _11019_ (.A(_01811_),
    .B(_01813_),
    .X(_01814_));
 sky130_fd_sc_hd__xnor2_4 _11020_ (.A(_01811_),
    .B(_01813_),
    .Y(_01815_));
 sky130_fd_sc_hd__or2_2 _11021_ (.A(_01806_),
    .B(_01815_),
    .X(_01816_));
 sky130_fd_sc_hd__xor2_4 _11022_ (.A(_01806_),
    .B(_01815_),
    .X(_01817_));
 sky130_fd_sc_hd__o21ai_4 _11023_ (.A1(_01763_),
    .A2(_01770_),
    .B1(_01817_),
    .Y(_01818_));
 sky130_fd_sc_hd__or3_2 _11024_ (.A(_01763_),
    .B(_01770_),
    .C(_01817_),
    .X(_01819_));
 sky130_fd_sc_hd__xnor2_1 _11025_ (.A(_01804_),
    .B(_01805_),
    .Y(_01820_));
 sky130_fd_sc_hd__nand2_4 _11026_ (.A(net447),
    .B(net913),
    .Y(_01821_));
 sky130_fd_sc_hd__and4_4 _11027_ (.A(net439),
    .B(net448),
    .C(net903),
    .D(net913),
    .X(_01822_));
 sky130_fd_sc_hd__a22oi_2 _11028_ (.A1(net447),
    .A2(net903),
    .B1(net918),
    .B2(net439),
    .Y(_01823_));
 sky130_fd_sc_hd__or3b_4 _11029_ (.A(_01822_),
    .B(_01823_),
    .C_N(_01820_),
    .X(_01824_));
 sky130_fd_sc_hd__xnor2_4 _11030_ (.A(_01498_),
    .B(_01500_),
    .Y(_01825_));
 sky130_fd_sc_hd__and2_2 _11031_ (.A(_01822_),
    .B(_01825_),
    .X(_01826_));
 sky130_fd_sc_hd__xnor2_4 _11032_ (.A(_01822_),
    .B(_01825_),
    .Y(_01827_));
 sky130_fd_sc_hd__a32o_4 _11033_ (.A1(net476),
    .A2(net873),
    .A3(_01802_),
    .B1(_01801_),
    .B2(net883),
    .X(_01828_));
 sky130_fd_sc_hd__and2b_2 _11034_ (.A_N(_01827_),
    .B(_01828_),
    .X(_01829_));
 sky130_fd_sc_hd__xor2_4 _11035_ (.A(_01827_),
    .B(_01828_),
    .X(_01830_));
 sky130_fd_sc_hd__xnor2_4 _11036_ (.A(_01490_),
    .B(_01492_),
    .Y(_01831_));
 sky130_fd_sc_hd__and2b_4 _11037_ (.A_N(_01830_),
    .B(_01831_),
    .X(_01832_));
 sky130_fd_sc_hd__xnor2_4 _11038_ (.A(_01830_),
    .B(_01831_),
    .Y(_01833_));
 sky130_fd_sc_hd__nand2b_2 _11039_ (.A_N(_01824_),
    .B(_01833_),
    .Y(_01834_));
 sky130_fd_sc_hd__xnor2_4 _11040_ (.A(_01824_),
    .B(_01833_),
    .Y(_01835_));
 sky130_fd_sc_hd__nand3_4 _11041_ (.A(_01818_),
    .B(_01819_),
    .C(_01835_),
    .Y(_01836_));
 sky130_fd_sc_hd__a21o_1 _11042_ (.A1(_01818_),
    .A2(_01819_),
    .B1(_01835_),
    .X(_01837_));
 sky130_fd_sc_hd__xnor2_4 _11043_ (.A(_01754_),
    .B(_01755_),
    .Y(_01838_));
 sky130_fd_sc_hd__nand2b_2 _11044_ (.A_N(_01821_),
    .B(_01838_),
    .Y(_01839_));
 sky130_fd_sc_hd__o21bai_1 _11045_ (.A1(_01822_),
    .A2(_01823_),
    .B1_N(_01820_),
    .Y(_01840_));
 sky130_fd_sc_hd__nand2_2 _11046_ (.A(_01824_),
    .B(_01840_),
    .Y(_01841_));
 sky130_fd_sc_hd__nor2_2 _11047_ (.A(_01839_),
    .B(_01841_),
    .Y(_01842_));
 sky130_fd_sc_hd__xor2_2 _11048_ (.A(_01839_),
    .B(_01841_),
    .X(_01843_));
 sky130_fd_sc_hd__or3_2 _11049_ (.A(_01712_),
    .B(_01720_),
    .C(_01773_),
    .X(_01844_));
 sky130_fd_sc_hd__and3_2 _11050_ (.A(_01774_),
    .B(_01843_),
    .C(_01844_),
    .X(_01845_));
 sky130_fd_sc_hd__nand3_2 _11051_ (.A(_01774_),
    .B(_01843_),
    .C(_01844_),
    .Y(_01846_));
 sky130_fd_sc_hd__o211ai_4 _11052_ (.A1(_01842_),
    .A2(_01845_),
    .B1(_01836_),
    .C1(_01837_),
    .Y(_01847_));
 sky130_fd_sc_hd__inv_2 _11053_ (.A(_01847_),
    .Y(_01848_));
 sky130_fd_sc_hd__a211o_2 _11054_ (.A1(_01836_),
    .A2(_01837_),
    .B1(_01842_),
    .C1(_01845_),
    .X(_01849_));
 sky130_fd_sc_hd__and4_4 _11055_ (.A(_01798_),
    .B(_01799_),
    .C(_01847_),
    .D(_01849_),
    .X(_01850_));
 sky130_fd_sc_hd__a22oi_4 _11056_ (.A1(_01798_),
    .A2(_01799_),
    .B1(_01847_),
    .B2(_01849_),
    .Y(_01851_));
 sky130_fd_sc_hd__nand3_2 _11057_ (.A(_01608_),
    .B(_01610_),
    .C(_01723_),
    .Y(_01852_));
 sky130_fd_sc_hd__xnor2_4 _11058_ (.A(_01821_),
    .B(_01838_),
    .Y(_01853_));
 sky130_fd_sc_hd__and3_4 _11059_ (.A(_01724_),
    .B(_01852_),
    .C(_01853_),
    .X(_01854_));
 sky130_fd_sc_hd__a21o_1 _11060_ (.A1(_01774_),
    .A2(_01844_),
    .B1(_01843_),
    .X(_01855_));
 sky130_fd_sc_hd__nand3_4 _11061_ (.A(_01846_),
    .B(_01854_),
    .C(_01855_),
    .Y(_01856_));
 sky130_fd_sc_hd__a211o_4 _11062_ (.A1(_01743_),
    .A2(_01744_),
    .B1(_01652_),
    .C1(_01656_),
    .X(_01857_));
 sky130_fd_sc_hd__a21o_2 _11063_ (.A1(_01846_),
    .A2(_01855_),
    .B1(_01854_),
    .X(_01858_));
 sky130_fd_sc_hd__and4_2 _11064_ (.A(_01745_),
    .B(_01856_),
    .C(_01857_),
    .D(_01858_),
    .X(_01859_));
 sky130_fd_sc_hd__nand4_4 _11065_ (.A(_01745_),
    .B(_01856_),
    .C(_01857_),
    .D(_01858_),
    .Y(_01860_));
 sky130_fd_sc_hd__a211oi_4 _11066_ (.A1(_01856_),
    .A2(_01860_),
    .B1(_01850_),
    .C1(_01851_),
    .Y(_01861_));
 sky130_fd_sc_hd__inv_2 _11067_ (.A(_01861_),
    .Y(_01862_));
 sky130_fd_sc_hd__o211a_2 _11068_ (.A1(_01850_),
    .A2(_01851_),
    .B1(_01856_),
    .C1(_01860_),
    .X(_01863_));
 sky130_fd_sc_hd__or3_4 _11069_ (.A(_01748_),
    .B(_01861_),
    .C(_01863_),
    .X(_01864_));
 sky130_fd_sc_hd__o21ai_4 _11070_ (.A1(_01861_),
    .A2(_01863_),
    .B1(_01748_),
    .Y(_01865_));
 sky130_fd_sc_hd__a22oi_4 _11071_ (.A1(_01745_),
    .A2(_01857_),
    .B1(_01858_),
    .B2(_01856_),
    .Y(_01866_));
 sky130_fd_sc_hd__and3_2 _11072_ (.A(_01611_),
    .B(_01618_),
    .C(_01625_),
    .X(_01867_));
 sky130_fd_sc_hd__or2_1 _11073_ (.A(_01699_),
    .B(_01704_),
    .X(_01868_));
 sky130_fd_sc_hd__nand2_2 _11074_ (.A(_01705_),
    .B(_01868_),
    .Y(_01869_));
 sky130_fd_sc_hd__or3_4 _11075_ (.A(_01627_),
    .B(_01867_),
    .C(_01869_),
    .X(_01870_));
 sky130_fd_sc_hd__a21oi_4 _11076_ (.A1(_01724_),
    .A2(_01852_),
    .B1(_01853_),
    .Y(_01871_));
 sky130_fd_sc_hd__or3_4 _11077_ (.A(_01854_),
    .B(_01870_),
    .C(_01871_),
    .X(_01872_));
 sky130_fd_sc_hd__a211o_2 _11078_ (.A1(_01658_),
    .A2(_01659_),
    .B1(_01676_),
    .C1(_01688_),
    .X(_01873_));
 sky130_fd_sc_hd__o21ai_4 _11079_ (.A1(_01854_),
    .A2(_01871_),
    .B1(_01870_),
    .Y(_01874_));
 sky130_fd_sc_hd__nand4_4 _11080_ (.A(_01689_),
    .B(_01872_),
    .C(_01873_),
    .D(_01874_),
    .Y(_01875_));
 sky130_fd_sc_hd__a211oi_4 _11081_ (.A1(_01872_),
    .A2(_01875_),
    .B1(_01859_),
    .C1(_01866_),
    .Y(_01876_));
 sky130_fd_sc_hd__xnor2_4 _11082_ (.A(_01591_),
    .B(_01690_),
    .Y(_01877_));
 sky130_fd_sc_hd__o211a_2 _11083_ (.A1(_01859_),
    .A2(_01866_),
    .B1(_01872_),
    .C1(_01875_),
    .X(_01878_));
 sky130_fd_sc_hd__nor3_4 _11084_ (.A(_01876_),
    .B(_01877_),
    .C(_01878_),
    .Y(_01879_));
 sky130_fd_sc_hd__o211a_1 _11085_ (.A1(_01876_),
    .A2(_01879_),
    .B1(_01864_),
    .C1(_01865_),
    .X(_01880_));
 sky130_fd_sc_hd__a211oi_4 _11086_ (.A1(_01864_),
    .A2(_01865_),
    .B1(_01876_),
    .C1(_01879_),
    .Y(_01881_));
 sky130_fd_sc_hd__nor2_2 _11087_ (.A(_01880_),
    .B(_01881_),
    .Y(_01882_));
 sky130_fd_sc_hd__xnor2_4 _11088_ (.A(_01691_),
    .B(_01882_),
    .Y(_01883_));
 sky130_fd_sc_hd__o21a_1 _11089_ (.A1(_01876_),
    .A2(_01878_),
    .B1(_01877_),
    .X(_01884_));
 sky130_fd_sc_hd__nor2_2 _11090_ (.A(_01879_),
    .B(_01884_),
    .Y(_01885_));
 sky130_fd_sc_hd__a22o_2 _11091_ (.A1(_01689_),
    .A2(_01873_),
    .B1(_01874_),
    .B2(_01872_),
    .X(_01886_));
 sky130_fd_sc_hd__xnor2_2 _11092_ (.A(_01623_),
    .B(_01624_),
    .Y(_01887_));
 sky130_fd_sc_hd__o2bb2a_1 _11093_ (.A1_N(net505),
    .A2_N(net888),
    .B1(_01614_),
    .B2(_01615_),
    .X(_01888_));
 sky130_fd_sc_hd__nor2_2 _11094_ (.A(_01616_),
    .B(_01888_),
    .Y(_01889_));
 sky130_fd_sc_hd__and4_2 _11095_ (.A(net488),
    .B(net498),
    .C(net908),
    .D(net916),
    .X(_01890_));
 sky130_fd_sc_hd__a22oi_2 _11096_ (.A1(net498),
    .A2(net908),
    .B1(net916),
    .B2(net488),
    .Y(_01891_));
 sky130_fd_sc_hd__and4bb_4 _11097_ (.A_N(_01890_),
    .B_N(_01891_),
    .C(net505),
    .D(net897),
    .X(_01892_));
 sky130_fd_sc_hd__nor2_4 _11098_ (.A(_01890_),
    .B(_01892_),
    .Y(_01893_));
 sky130_fd_sc_hd__or3_2 _11099_ (.A(_01616_),
    .B(_01888_),
    .C(_01893_),
    .X(_01894_));
 sky130_fd_sc_hd__xnor2_4 _11100_ (.A(_01663_),
    .B(_01665_),
    .Y(_01895_));
 sky130_fd_sc_hd__xnor2_4 _11101_ (.A(_01889_),
    .B(_01893_),
    .Y(_01896_));
 sky130_fd_sc_hd__nand2_1 _11102_ (.A(_01895_),
    .B(_01896_),
    .Y(_01897_));
 sky130_fd_sc_hd__a21o_2 _11103_ (.A1(_01894_),
    .A2(_01897_),
    .B1(_01887_),
    .X(_01898_));
 sky130_fd_sc_hd__nand3_2 _11104_ (.A(_01887_),
    .B(_01894_),
    .C(_01897_),
    .Y(_01899_));
 sky130_fd_sc_hd__nand2_4 _11105_ (.A(_01898_),
    .B(_01899_),
    .Y(_01900_));
 sky130_fd_sc_hd__a22oi_1 _11106_ (.A1(net475),
    .A2(net903),
    .B1(net913),
    .B2(net466),
    .Y(_01901_));
 sky130_fd_sc_hd__or2_4 _11107_ (.A(_01699_),
    .B(_01901_),
    .X(_01902_));
 sky130_fd_sc_hd__nor2_2 _11108_ (.A(_01900_),
    .B(_01902_),
    .Y(_01903_));
 sky130_fd_sc_hd__o21ai_4 _11109_ (.A1(_01627_),
    .A2(_01867_),
    .B1(_01869_),
    .Y(_01904_));
 sky130_fd_sc_hd__nand3_4 _11110_ (.A(_01870_),
    .B(_01903_),
    .C(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__a21oi_4 _11111_ (.A1(_01677_),
    .A2(_01678_),
    .B1(_01687_),
    .Y(_01906_));
 sky130_fd_sc_hd__or3_4 _11112_ (.A(_01688_),
    .B(_01898_),
    .C(_01906_),
    .X(_01907_));
 sky130_fd_sc_hd__o21ai_4 _11113_ (.A1(_01688_),
    .A2(_01906_),
    .B1(_01898_),
    .Y(_01908_));
 sky130_fd_sc_hd__xnor2_4 _11114_ (.A(_01673_),
    .B(_01674_),
    .Y(_01909_));
 sky130_fd_sc_hd__and4_2 _11115_ (.A(net512),
    .B(net524),
    .C(net877),
    .D(net888),
    .X(_01910_));
 sky130_fd_sc_hd__a22oi_2 _11116_ (.A1(net524),
    .A2(net877),
    .B1(net888),
    .B2(net512),
    .Y(_01911_));
 sky130_fd_sc_hd__and4bb_4 _11117_ (.A_N(_01910_),
    .B_N(_01911_),
    .C(net529),
    .D(net866),
    .X(_01912_));
 sky130_fd_sc_hd__nor2_4 _11118_ (.A(_01910_),
    .B(_01912_),
    .Y(_01913_));
 sky130_fd_sc_hd__o2bb2a_1 _11119_ (.A1_N(net573),
    .A2_N(net825),
    .B1(_01670_),
    .B2(_01671_),
    .X(_01914_));
 sky130_fd_sc_hd__nor2_2 _11120_ (.A(_01672_),
    .B(_01914_),
    .Y(_01915_));
 sky130_fd_sc_hd__or3_4 _11121_ (.A(_01672_),
    .B(_01913_),
    .C(_01914_),
    .X(_01916_));
 sky130_fd_sc_hd__and4_1 _11122_ (.A(net542),
    .B(net556),
    .C(net846),
    .D(net856),
    .X(_01917_));
 sky130_fd_sc_hd__a22oi_2 _11123_ (.A1(net556),
    .A2(net846),
    .B1(net856),
    .B2(net542),
    .Y(_01918_));
 sky130_fd_sc_hd__and4bb_2 _11124_ (.A_N(_01917_),
    .B_N(_01918_),
    .C(net573),
    .D(net835),
    .X(_01919_));
 sky130_fd_sc_hd__or2_4 _11125_ (.A(_01917_),
    .B(_01919_),
    .X(_01920_));
 sky130_fd_sc_hd__xnor2_4 _11126_ (.A(_01913_),
    .B(_01915_),
    .Y(_01921_));
 sky130_fd_sc_hd__nand2_2 _11127_ (.A(_01920_),
    .B(_01921_),
    .Y(_01922_));
 sky130_fd_sc_hd__a21oi_4 _11128_ (.A1(_01916_),
    .A2(_01922_),
    .B1(_01909_),
    .Y(_01923_));
 sky130_fd_sc_hd__a21o_1 _11129_ (.A1(_01916_),
    .A2(_01922_),
    .B1(_01909_),
    .X(_01924_));
 sky130_fd_sc_hd__nand3_2 _11130_ (.A(_01909_),
    .B(_01916_),
    .C(_01922_),
    .Y(_01925_));
 sky130_fd_sc_hd__xnor2_4 _11131_ (.A(_01681_),
    .B(_01683_),
    .Y(_01926_));
 sky130_fd_sc_hd__and4_2 _11132_ (.A(net589),
    .B(net613),
    .C(net792),
    .D(net816),
    .X(_01927_));
 sky130_fd_sc_hd__a22oi_1 _11133_ (.A1(net613),
    .A2(net792),
    .B1(net817),
    .B2(net589),
    .Y(_01928_));
 sky130_fd_sc_hd__nor2_1 _11134_ (.A(_01927_),
    .B(_01928_),
    .Y(_01929_));
 sky130_fd_sc_hd__and3_2 _11135_ (.A(net602),
    .B(net805),
    .C(_01929_),
    .X(_01930_));
 sky130_fd_sc_hd__o21ai_4 _11136_ (.A1(_01927_),
    .A2(_01930_),
    .B1(_01926_),
    .Y(_01931_));
 sky130_fd_sc_hd__or3_1 _11137_ (.A(_01926_),
    .B(_01927_),
    .C(_01930_),
    .X(_01932_));
 sky130_fd_sc_hd__and2_2 _11138_ (.A(_01931_),
    .B(_01932_),
    .X(_01933_));
 sky130_fd_sc_hd__and3_4 _11139_ (.A(_01924_),
    .B(_01925_),
    .C(_01933_),
    .X(_01934_));
 sky130_fd_sc_hd__o211ai_4 _11140_ (.A1(_01923_),
    .A2(_01934_),
    .B1(_01907_),
    .C1(_01908_),
    .Y(_01935_));
 sky130_fd_sc_hd__a211o_2 _11141_ (.A1(_01907_),
    .A2(_01908_),
    .B1(_01923_),
    .C1(_01934_),
    .X(_01936_));
 sky130_fd_sc_hd__a21o_1 _11142_ (.A1(_01870_),
    .A2(_01904_),
    .B1(_01903_),
    .X(_01937_));
 sky130_fd_sc_hd__nand4_4 _11143_ (.A(_01905_),
    .B(_01935_),
    .C(_01936_),
    .D(_01937_),
    .Y(_01938_));
 sky130_fd_sc_hd__nand2_2 _11144_ (.A(_01905_),
    .B(_01938_),
    .Y(_01939_));
 sky130_fd_sc_hd__and3_4 _11145_ (.A(_01875_),
    .B(_01886_),
    .C(_01939_),
    .X(_01940_));
 sky130_fd_sc_hd__and2_1 _11146_ (.A(_01907_),
    .B(_01935_),
    .X(_01941_));
 sky130_fd_sc_hd__or2_4 _11147_ (.A(_01685_),
    .B(_01941_),
    .X(_01942_));
 sky130_fd_sc_hd__nand2_1 _11148_ (.A(_01685_),
    .B(_01941_),
    .Y(_01943_));
 sky130_fd_sc_hd__nand2_2 _11149_ (.A(_01942_),
    .B(_01943_),
    .Y(_01944_));
 sky130_fd_sc_hd__a21oi_4 _11150_ (.A1(_01875_),
    .A2(_01886_),
    .B1(_01939_),
    .Y(_01945_));
 sky130_fd_sc_hd__nor3_4 _11151_ (.A(_01940_),
    .B(_01944_),
    .C(_01945_),
    .Y(_01946_));
 sky130_fd_sc_hd__o21a_4 _11152_ (.A1(_01940_),
    .A2(_01946_),
    .B1(_01885_),
    .X(_01947_));
 sky130_fd_sc_hd__nor3_2 _11153_ (.A(_01885_),
    .B(_01940_),
    .C(_01946_),
    .Y(_01948_));
 sky130_fd_sc_hd__nor3_4 _11154_ (.A(_01942_),
    .B(_01947_),
    .C(_01948_),
    .Y(_01949_));
 sky130_fd_sc_hd__nor2_2 _11155_ (.A(_01947_),
    .B(_01949_),
    .Y(_01950_));
 sky130_fd_sc_hd__o21ai_4 _11156_ (.A1(_01947_),
    .A2(_01949_),
    .B1(_01883_),
    .Y(_01951_));
 sky130_fd_sc_hd__and2_2 _11157_ (.A(_01796_),
    .B(_01798_),
    .X(_01952_));
 sky130_fd_sc_hd__or2_4 _11158_ (.A(_01791_),
    .B(_01952_),
    .X(_01953_));
 sky130_fd_sc_hd__xnor2_4 _11159_ (.A(_01791_),
    .B(_01952_),
    .Y(_01954_));
 sky130_fd_sc_hd__xnor2_2 _11160_ (.A(_01541_),
    .B(_01542_),
    .Y(_01955_));
 sky130_fd_sc_hd__a21oi_4 _11161_ (.A1(_01779_),
    .A2(_01781_),
    .B1(_01955_),
    .Y(_01956_));
 sky130_fd_sc_hd__and3_2 _11162_ (.A(_01779_),
    .B(_01781_),
    .C(_01955_),
    .X(_01957_));
 sky130_fd_sc_hd__o2bb2a_1 _11163_ (.A1_N(net599),
    .A2_N(net741),
    .B1(_01548_),
    .B2(_01549_),
    .X(_01958_));
 sky130_fd_sc_hd__nor2_1 _11164_ (.A(_01786_),
    .B(_01788_),
    .Y(_01959_));
 sky130_fd_sc_hd__or3_1 _11165_ (.A(_01550_),
    .B(_01958_),
    .C(_01959_),
    .X(_01960_));
 sky130_fd_sc_hd__o21ai_1 _11166_ (.A1(_01550_),
    .A2(_01958_),
    .B1(_01959_),
    .Y(_01961_));
 sky130_fd_sc_hd__and2_1 _11167_ (.A(_01960_),
    .B(_01961_),
    .X(_01962_));
 sky130_fd_sc_hd__nor3b_4 _11168_ (.A(_01956_),
    .B(_01957_),
    .C_N(_01962_),
    .Y(_01963_));
 sky130_fd_sc_hd__o21ba_2 _11169_ (.A1(_01956_),
    .A2(_01957_),
    .B1_N(_01962_),
    .X(_01964_));
 sky130_fd_sc_hd__a211o_2 _11170_ (.A1(_01816_),
    .A2(_01818_),
    .B1(_01963_),
    .C1(_01964_),
    .X(_01965_));
 sky130_fd_sc_hd__o211ai_4 _11171_ (.A1(_01963_),
    .A2(_01964_),
    .B1(_01816_),
    .C1(_01818_),
    .Y(_01966_));
 sky130_fd_sc_hd__o211ai_4 _11172_ (.A1(_01783_),
    .A2(_01794_),
    .B1(_01965_),
    .C1(_01966_),
    .Y(_01967_));
 sky130_fd_sc_hd__a211o_2 _11173_ (.A1(_01965_),
    .A2(_01966_),
    .B1(_01783_),
    .C1(_01794_),
    .X(_01968_));
 sky130_fd_sc_hd__xor2_4 _11174_ (.A(_01517_),
    .B(_01519_),
    .X(_01969_));
 sky130_fd_sc_hd__o21ai_4 _11175_ (.A1(_01826_),
    .A2(_01829_),
    .B1(_01969_),
    .Y(_01970_));
 sky130_fd_sc_hd__or3_4 _11176_ (.A(_01826_),
    .B(_01829_),
    .C(_01969_),
    .X(_01971_));
 sky130_fd_sc_hd__o211a_2 _11177_ (.A1(_01810_),
    .A2(_01814_),
    .B1(_01970_),
    .C1(_01971_),
    .X(_01972_));
 sky130_fd_sc_hd__o211ai_4 _11178_ (.A1(_01810_),
    .A2(_01814_),
    .B1(_01970_),
    .C1(_01971_),
    .Y(_01973_));
 sky130_fd_sc_hd__a211oi_4 _11179_ (.A1(_01970_),
    .A2(_01971_),
    .B1(_01810_),
    .C1(_01814_),
    .Y(_01974_));
 sky130_fd_sc_hd__xor2_4 _11180_ (.A(_01503_),
    .B(_01504_),
    .X(_01975_));
 sky130_fd_sc_hd__xnor2_4 _11181_ (.A(_01832_),
    .B(_01975_),
    .Y(_01976_));
 sky130_fd_sc_hd__nor3_4 _11182_ (.A(_01972_),
    .B(_01974_),
    .C(_01976_),
    .Y(_01977_));
 sky130_fd_sc_hd__o21a_2 _11183_ (.A1(_01972_),
    .A2(_01974_),
    .B1(_01976_),
    .X(_01978_));
 sky130_fd_sc_hd__a211o_4 _11184_ (.A1(_01834_),
    .A2(_01836_),
    .B1(_01977_),
    .C1(_01978_),
    .X(_01979_));
 sky130_fd_sc_hd__o211ai_4 _11185_ (.A1(_01977_),
    .A2(_01978_),
    .B1(_01834_),
    .C1(_01836_),
    .Y(_01980_));
 sky130_fd_sc_hd__nand4_4 _11186_ (.A(_01967_),
    .B(_01968_),
    .C(_01979_),
    .D(_01980_),
    .Y(_01981_));
 sky130_fd_sc_hd__a22o_2 _11187_ (.A1(_01967_),
    .A2(_01968_),
    .B1(_01979_),
    .B2(_01980_),
    .X(_01982_));
 sky130_fd_sc_hd__o211a_2 _11188_ (.A1(_01848_),
    .A2(_01850_),
    .B1(_01981_),
    .C1(_01982_),
    .X(_01983_));
 sky130_fd_sc_hd__a211oi_4 _11189_ (.A1(_01981_),
    .A2(_01982_),
    .B1(_01848_),
    .C1(_01850_),
    .Y(_01984_));
 sky130_fd_sc_hd__nor3_4 _11190_ (.A(_01954_),
    .B(_01983_),
    .C(_01984_),
    .Y(_01985_));
 sky130_fd_sc_hd__o21a_2 _11191_ (.A1(_01983_),
    .A2(_01984_),
    .B1(_01954_),
    .X(_01986_));
 sky130_fd_sc_hd__a211oi_4 _11192_ (.A1(_01862_),
    .A2(_01864_),
    .B1(_01985_),
    .C1(_01986_),
    .Y(_01987_));
 sky130_fd_sc_hd__o211a_2 _11193_ (.A1(_01985_),
    .A2(_01986_),
    .B1(_01862_),
    .C1(_01864_),
    .X(_01988_));
 sky130_fd_sc_hd__nor2_2 _11194_ (.A(_01987_),
    .B(_01988_),
    .Y(_01989_));
 sky130_fd_sc_hd__xnor2_4 _11195_ (.A(_01747_),
    .B(_01989_),
    .Y(_01990_));
 sky130_fd_sc_hd__o21ba_2 _11196_ (.A1(_01691_),
    .A2(_01881_),
    .B1_N(_01880_),
    .X(_01991_));
 sky130_fd_sc_hd__and2b_2 _11197_ (.A_N(_01991_),
    .B(_01990_),
    .X(_01992_));
 sky130_fd_sc_hd__xnor2_4 _11198_ (.A(_01990_),
    .B(_01991_),
    .Y(_01993_));
 sky130_fd_sc_hd__and2b_1 _11199_ (.A_N(_01951_),
    .B(_01993_),
    .X(_01994_));
 sky130_fd_sc_hd__nand2b_1 _11200_ (.A_N(_01951_),
    .B(_01993_),
    .Y(_01995_));
 sky130_fd_sc_hd__xnor2_4 _11201_ (.A(_01951_),
    .B(_01993_),
    .Y(_01996_));
 sky130_fd_sc_hd__and2_1 _11202_ (.A(_01965_),
    .B(_01967_),
    .X(_01997_));
 sky130_fd_sc_hd__or2_2 _11203_ (.A(_01960_),
    .B(_01997_),
    .X(_01998_));
 sky130_fd_sc_hd__nand2_1 _11204_ (.A(_01960_),
    .B(_01997_),
    .Y(_01999_));
 sky130_fd_sc_hd__nand2_4 _11205_ (.A(_01998_),
    .B(_01999_),
    .Y(_02000_));
 sky130_fd_sc_hd__a21oi_4 _11206_ (.A1(_01544_),
    .A2(_01545_),
    .B1(_01554_),
    .Y(_02001_));
 sky130_fd_sc_hd__a211o_2 _11207_ (.A1(_01970_),
    .A2(_01973_),
    .B1(_02001_),
    .C1(_01555_),
    .X(_02002_));
 sky130_fd_sc_hd__o211ai_4 _11208_ (.A1(_01555_),
    .A2(_02001_),
    .B1(_01973_),
    .C1(_01970_),
    .Y(_02003_));
 sky130_fd_sc_hd__o211ai_4 _11209_ (.A1(_01956_),
    .A2(_01963_),
    .B1(_02002_),
    .C1(_02003_),
    .Y(_02004_));
 sky130_fd_sc_hd__a211o_1 _11210_ (.A1(_02002_),
    .A2(_02003_),
    .B1(_01956_),
    .C1(_01963_),
    .X(_02005_));
 sky130_fd_sc_hd__nand2_4 _11211_ (.A(_02004_),
    .B(_02005_),
    .Y(_02006_));
 sky130_fd_sc_hd__xnor2_4 _11212_ (.A(_01523_),
    .B(_01524_),
    .Y(_02007_));
 sky130_fd_sc_hd__a21o_2 _11213_ (.A1(_01832_),
    .A2(_01975_),
    .B1(_01977_),
    .X(_02008_));
 sky130_fd_sc_hd__nand2_1 _11214_ (.A(_02007_),
    .B(_02008_),
    .Y(_02009_));
 sky130_fd_sc_hd__nor2_1 _11215_ (.A(_02007_),
    .B(_02008_),
    .Y(_02010_));
 sky130_fd_sc_hd__xor2_4 _11216_ (.A(_02007_),
    .B(_02008_),
    .X(_02011_));
 sky130_fd_sc_hd__xnor2_4 _11217_ (.A(_02006_),
    .B(_02011_),
    .Y(_02012_));
 sky130_fd_sc_hd__nand2_4 _11218_ (.A(_01979_),
    .B(_01981_),
    .Y(_02013_));
 sky130_fd_sc_hd__nand2_1 _11219_ (.A(_02012_),
    .B(_02013_),
    .Y(_02014_));
 sky130_fd_sc_hd__xnor2_4 _11220_ (.A(_02012_),
    .B(_02013_),
    .Y(_02015_));
 sky130_fd_sc_hd__xor2_4 _11221_ (.A(_02000_),
    .B(_02015_),
    .X(_02016_));
 sky130_fd_sc_hd__or2_4 _11222_ (.A(_01983_),
    .B(_01985_),
    .X(_02017_));
 sky130_fd_sc_hd__xor2_4 _11223_ (.A(_02016_),
    .B(_02017_),
    .X(_02018_));
 sky130_fd_sc_hd__and2b_1 _11224_ (.A_N(_01953_),
    .B(_02018_),
    .X(_02019_));
 sky130_fd_sc_hd__xnor2_4 _11225_ (.A(_01953_),
    .B(_02018_),
    .Y(_02020_));
 sky130_fd_sc_hd__o21bai_4 _11226_ (.A1(_01747_),
    .A2(_01988_),
    .B1_N(_01987_),
    .Y(_02021_));
 sky130_fd_sc_hd__and2_4 _11227_ (.A(_02020_),
    .B(_02021_),
    .X(_02022_));
 sky130_fd_sc_hd__xor2_4 _11228_ (.A(_02020_),
    .B(_02021_),
    .X(_02023_));
 sky130_fd_sc_hd__xnor2_2 _11229_ (.A(_01992_),
    .B(_02023_),
    .Y(_02024_));
 sky130_fd_sc_hd__and2b_1 _11230_ (.A_N(_02024_),
    .B(_01996_),
    .X(_02025_));
 sky130_fd_sc_hd__o21a_1 _11231_ (.A1(_01992_),
    .A2(_01994_),
    .B1(_02023_),
    .X(_02026_));
 sky130_fd_sc_hd__xnor2_4 _11232_ (.A(_01883_),
    .B(_01950_),
    .Y(_02027_));
 sky130_fd_sc_hd__o21a_1 _11233_ (.A1(_01947_),
    .A2(_01948_),
    .B1(_01942_),
    .X(_02028_));
 sky130_fd_sc_hd__or2_4 _11234_ (.A(_01949_),
    .B(_02028_),
    .X(_02029_));
 sky130_fd_sc_hd__o21a_2 _11235_ (.A1(_01940_),
    .A2(_01945_),
    .B1(_01944_),
    .X(_02030_));
 sky130_fd_sc_hd__a22o_1 _11236_ (.A1(_01935_),
    .A2(_01936_),
    .B1(_01937_),
    .B2(_01905_),
    .X(_02031_));
 sky130_fd_sc_hd__nand2_4 _11237_ (.A(_01938_),
    .B(_02031_),
    .Y(_02032_));
 sky130_fd_sc_hd__xor2_4 _11238_ (.A(_01895_),
    .B(_01896_),
    .X(_02033_));
 sky130_fd_sc_hd__nand2_4 _11239_ (.A(net507),
    .B(net916),
    .Y(_02034_));
 sky130_fd_sc_hd__and4_4 _11240_ (.A(net498),
    .B(net505),
    .C(net908),
    .D(net916),
    .X(_02035_));
 sky130_fd_sc_hd__o2bb2a_1 _11241_ (.A1_N(net505),
    .A2_N(net897),
    .B1(_01890_),
    .B2(_01891_),
    .X(_02036_));
 sky130_fd_sc_hd__nor2_4 _11242_ (.A(_01892_),
    .B(_02036_),
    .Y(_02037_));
 sky130_fd_sc_hd__and2_2 _11243_ (.A(_02035_),
    .B(_02037_),
    .X(_02038_));
 sky130_fd_sc_hd__xnor2_4 _11244_ (.A(_02035_),
    .B(_02037_),
    .Y(_02039_));
 sky130_fd_sc_hd__o2bb2a_1 _11245_ (.A1_N(net530),
    .A2_N(net866),
    .B1(_01910_),
    .B2(_01911_),
    .X(_02040_));
 sky130_fd_sc_hd__nor2_4 _11246_ (.A(_01912_),
    .B(_02040_),
    .Y(_02041_));
 sky130_fd_sc_hd__and2b_1 _11247_ (.A_N(_02039_),
    .B(_02041_),
    .X(_02042_));
 sky130_fd_sc_hd__o21ai_4 _11248_ (.A1(_02038_),
    .A2(_02042_),
    .B1(_02033_),
    .Y(_02043_));
 sky130_fd_sc_hd__or3_1 _11249_ (.A(_02033_),
    .B(_02038_),
    .C(_02042_),
    .X(_02044_));
 sky130_fd_sc_hd__nand2_1 _11250_ (.A(_02043_),
    .B(_02044_),
    .Y(_02045_));
 sky130_fd_sc_hd__or2_4 _11251_ (.A(_01698_),
    .B(_02045_),
    .X(_02046_));
 sky130_fd_sc_hd__xnor2_4 _11252_ (.A(_01900_),
    .B(_01902_),
    .Y(_02047_));
 sky130_fd_sc_hd__xor2_4 _11253_ (.A(_02046_),
    .B(_02047_),
    .X(_02048_));
 sky130_fd_sc_hd__a21oi_4 _11254_ (.A1(_01924_),
    .A2(_01925_),
    .B1(_01933_),
    .Y(_02049_));
 sky130_fd_sc_hd__or3_4 _11255_ (.A(_01934_),
    .B(_02043_),
    .C(_02049_),
    .X(_02050_));
 sky130_fd_sc_hd__o21ai_4 _11256_ (.A1(_01934_),
    .A2(_02049_),
    .B1(_02043_),
    .Y(_02051_));
 sky130_fd_sc_hd__xnor2_4 _11257_ (.A(_01920_),
    .B(_01921_),
    .Y(_02052_));
 sky130_fd_sc_hd__and4_2 _11258_ (.A(net515),
    .B(net522),
    .C(net888),
    .D(net897),
    .X(_02053_));
 sky130_fd_sc_hd__a22oi_2 _11259_ (.A1(net522),
    .A2(net888),
    .B1(net897),
    .B2(net515),
    .Y(_02054_));
 sky130_fd_sc_hd__and4bb_2 _11260_ (.A_N(_02053_),
    .B_N(_02054_),
    .C(net530),
    .D(net877),
    .X(_02055_));
 sky130_fd_sc_hd__nor2_4 _11261_ (.A(_02053_),
    .B(_02055_),
    .Y(_02056_));
 sky130_fd_sc_hd__o2bb2a_1 _11262_ (.A1_N(net573),
    .A2_N(net835),
    .B1(_01917_),
    .B2(_01918_),
    .X(_02057_));
 sky130_fd_sc_hd__nor2_2 _11263_ (.A(_01919_),
    .B(_02057_),
    .Y(_02058_));
 sky130_fd_sc_hd__or3_4 _11264_ (.A(_01919_),
    .B(_02056_),
    .C(_02057_),
    .X(_02059_));
 sky130_fd_sc_hd__and2_2 _11265_ (.A(net545),
    .B(net865),
    .X(_02060_));
 sky130_fd_sc_hd__nand4_4 _11266_ (.A(net546),
    .B(net561),
    .C(net856),
    .D(net866),
    .Y(_02061_));
 sky130_fd_sc_hd__a22o_2 _11267_ (.A1(net560),
    .A2(net856),
    .B1(net866),
    .B2(net546),
    .X(_02062_));
 sky130_fd_sc_hd__and4_2 _11268_ (.A(net579),
    .B(net846),
    .C(_02061_),
    .D(_02062_),
    .X(_02063_));
 sky130_fd_sc_hd__a31o_4 _11269_ (.A1(net560),
    .A2(net856),
    .A3(_02060_),
    .B1(_02063_),
    .X(_02064_));
 sky130_fd_sc_hd__xnor2_4 _11270_ (.A(_02056_),
    .B(_02058_),
    .Y(_02065_));
 sky130_fd_sc_hd__nand2_2 _11271_ (.A(_02064_),
    .B(_02065_),
    .Y(_02066_));
 sky130_fd_sc_hd__a21oi_4 _11272_ (.A1(_02059_),
    .A2(_02066_),
    .B1(_02052_),
    .Y(_02067_));
 sky130_fd_sc_hd__a21o_1 _11273_ (.A1(_02059_),
    .A2(_02066_),
    .B1(_02052_),
    .X(_02068_));
 sky130_fd_sc_hd__nand3_2 _11274_ (.A(_02052_),
    .B(_02059_),
    .C(_02066_),
    .Y(_02069_));
 sky130_fd_sc_hd__a21o_1 _11275_ (.A1(net602),
    .A2(net805),
    .B1(_01929_),
    .X(_02070_));
 sky130_fd_sc_hd__and2b_1 _11276_ (.A_N(_01930_),
    .B(_02070_),
    .X(_02071_));
 sky130_fd_sc_hd__and2_2 _11277_ (.A(net612),
    .B(net827),
    .X(_02072_));
 sky130_fd_sc_hd__and3_2 _11278_ (.A(net591),
    .B(net808),
    .C(_02072_),
    .X(_02073_));
 sky130_fd_sc_hd__a22oi_1 _11279_ (.A1(net613),
    .A2(net808),
    .B1(net827),
    .B2(net589),
    .Y(_02074_));
 sky130_fd_sc_hd__nor2_1 _11280_ (.A(_02073_),
    .B(_02074_),
    .Y(_02075_));
 sky130_fd_sc_hd__and3_4 _11281_ (.A(net604),
    .B(net817),
    .C(_02075_),
    .X(_02076_));
 sky130_fd_sc_hd__o21ai_4 _11282_ (.A1(_02073_),
    .A2(_02076_),
    .B1(_02071_),
    .Y(_02077_));
 sky130_fd_sc_hd__or3_1 _11283_ (.A(_02071_),
    .B(_02073_),
    .C(_02076_),
    .X(_02078_));
 sky130_fd_sc_hd__and2_2 _11284_ (.A(_02077_),
    .B(_02078_),
    .X(_02079_));
 sky130_fd_sc_hd__and3_4 _11285_ (.A(_02068_),
    .B(_02069_),
    .C(_02079_),
    .X(_02080_));
 sky130_fd_sc_hd__o211ai_4 _11286_ (.A1(_02067_),
    .A2(_02080_),
    .B1(_02050_),
    .C1(_02051_),
    .Y(_02081_));
 sky130_fd_sc_hd__a211o_2 _11287_ (.A1(_02050_),
    .A2(_02051_),
    .B1(_02067_),
    .C1(_02080_),
    .X(_02082_));
 sky130_fd_sc_hd__nand3_4 _11288_ (.A(_02048_),
    .B(_02081_),
    .C(_02082_),
    .Y(_02083_));
 sky130_fd_sc_hd__o21ai_4 _11289_ (.A1(_02046_),
    .A2(_02047_),
    .B1(_02083_),
    .Y(_02084_));
 sky130_fd_sc_hd__nand2b_2 _11290_ (.A_N(_02032_),
    .B(_02084_),
    .Y(_02085_));
 sky130_fd_sc_hd__and2_1 _11291_ (.A(_02050_),
    .B(_02081_),
    .X(_02086_));
 sky130_fd_sc_hd__or2_4 _11292_ (.A(_01931_),
    .B(_02086_),
    .X(_02087_));
 sky130_fd_sc_hd__nand2_1 _11293_ (.A(_01931_),
    .B(_02086_),
    .Y(_02088_));
 sky130_fd_sc_hd__nand2_4 _11294_ (.A(_02087_),
    .B(_02088_),
    .Y(_02089_));
 sky130_fd_sc_hd__xnor2_4 _11295_ (.A(_02032_),
    .B(_02084_),
    .Y(_02090_));
 sky130_fd_sc_hd__nand2b_2 _11296_ (.A_N(_02089_),
    .B(_02090_),
    .Y(_02091_));
 sky130_fd_sc_hd__a211oi_4 _11297_ (.A1(_02085_),
    .A2(_02091_),
    .B1(_01946_),
    .C1(_02030_),
    .Y(_02092_));
 sky130_fd_sc_hd__o211a_1 _11298_ (.A1(_01946_),
    .A2(_02030_),
    .B1(_02085_),
    .C1(_02091_),
    .X(_02093_));
 sky130_fd_sc_hd__or3_4 _11299_ (.A(_02087_),
    .B(_02092_),
    .C(_02093_),
    .X(_02094_));
 sky130_fd_sc_hd__nand2b_4 _11300_ (.A_N(_02092_),
    .B(_02094_),
    .Y(_02095_));
 sky130_fd_sc_hd__and2b_2 _11301_ (.A_N(_02029_),
    .B(_02095_),
    .X(_02096_));
 sky130_fd_sc_hd__xor2_4 _11302_ (.A(_02027_),
    .B(_02096_),
    .X(_02097_));
 sky130_fd_sc_hd__o2bb2a_1 _11303_ (.A1_N(net530),
    .A2_N(net877),
    .B1(_02053_),
    .B2(_02054_),
    .X(_02098_));
 sky130_fd_sc_hd__nor2_2 _11304_ (.A(_02055_),
    .B(_02098_),
    .Y(_02099_));
 sky130_fd_sc_hd__a22oi_2 _11305_ (.A1(net504),
    .A2(net908),
    .B1(net916),
    .B2(net498),
    .Y(_02100_));
 sky130_fd_sc_hd__nor2_2 _11306_ (.A(_02035_),
    .B(_02100_),
    .Y(_02101_));
 sky130_fd_sc_hd__nand2_4 _11307_ (.A(_02099_),
    .B(_02101_),
    .Y(_02102_));
 sky130_fd_sc_hd__xnor2_4 _11308_ (.A(_02039_),
    .B(_02041_),
    .Y(_02103_));
 sky130_fd_sc_hd__nand2b_2 _11309_ (.A_N(_02102_),
    .B(_02103_),
    .Y(_02104_));
 sky130_fd_sc_hd__a21oi_4 _11310_ (.A1(_02068_),
    .A2(_02069_),
    .B1(_02079_),
    .Y(_02105_));
 sky130_fd_sc_hd__or3_4 _11311_ (.A(_02080_),
    .B(_02104_),
    .C(_02105_),
    .X(_02106_));
 sky130_fd_sc_hd__o21ai_4 _11312_ (.A1(_02080_),
    .A2(_02105_),
    .B1(_02104_),
    .Y(_02107_));
 sky130_fd_sc_hd__xnor2_4 _11313_ (.A(_02064_),
    .B(_02065_),
    .Y(_02108_));
 sky130_fd_sc_hd__and4_1 _11314_ (.A(net515),
    .B(net522),
    .C(net897),
    .D(net907),
    .X(_02109_));
 sky130_fd_sc_hd__nand2_2 _11315_ (.A(net532),
    .B(net887),
    .Y(_02110_));
 sky130_fd_sc_hd__a22o_1 _11316_ (.A1(net522),
    .A2(net897),
    .B1(net907),
    .B2(net513),
    .X(_02111_));
 sky130_fd_sc_hd__and2b_2 _11317_ (.A_N(_02109_),
    .B(_02111_),
    .X(_02112_));
 sky130_fd_sc_hd__a31oi_2 _11318_ (.A1(net532),
    .A2(net887),
    .A3(_02111_),
    .B1(_02109_),
    .Y(_02113_));
 sky130_fd_sc_hd__a22oi_4 _11319_ (.A1(net578),
    .A2(net846),
    .B1(_02061_),
    .B2(_02062_),
    .Y(_02114_));
 sky130_fd_sc_hd__or3_4 _11320_ (.A(_02063_),
    .B(_02113_),
    .C(_02114_),
    .X(_02115_));
 sky130_fd_sc_hd__and2_1 _11321_ (.A(net560),
    .B(net876),
    .X(_02116_));
 sky130_fd_sc_hd__nand4_4 _11322_ (.A(net546),
    .B(net561),
    .C(net866),
    .D(net877),
    .Y(_02117_));
 sky130_fd_sc_hd__a22o_2 _11323_ (.A1(net561),
    .A2(net866),
    .B1(net877),
    .B2(net546),
    .X(_02118_));
 sky130_fd_sc_hd__nand4_4 _11324_ (.A(net578),
    .B(net856),
    .C(_02117_),
    .D(_02118_),
    .Y(_02119_));
 sky130_fd_sc_hd__nand2_4 _11325_ (.A(_02117_),
    .B(_02119_),
    .Y(_02120_));
 sky130_fd_sc_hd__o21ai_1 _11326_ (.A1(_02063_),
    .A2(_02114_),
    .B1(_02113_),
    .Y(_02121_));
 sky130_fd_sc_hd__and2_2 _11327_ (.A(_02115_),
    .B(_02121_),
    .X(_02122_));
 sky130_fd_sc_hd__nand2_2 _11328_ (.A(_02120_),
    .B(_02122_),
    .Y(_02123_));
 sky130_fd_sc_hd__a21oi_4 _11329_ (.A1(_02115_),
    .A2(_02123_),
    .B1(_02108_),
    .Y(_02124_));
 sky130_fd_sc_hd__a21o_1 _11330_ (.A1(_02115_),
    .A2(_02123_),
    .B1(_02108_),
    .X(_02125_));
 sky130_fd_sc_hd__nand3_2 _11331_ (.A(_02108_),
    .B(_02115_),
    .C(_02123_),
    .Y(_02126_));
 sky130_fd_sc_hd__a21oi_2 _11332_ (.A1(net604),
    .A2(net817),
    .B1(_02075_),
    .Y(_02127_));
 sky130_fd_sc_hd__nor2_4 _11333_ (.A(_02076_),
    .B(_02127_),
    .Y(_02128_));
 sky130_fd_sc_hd__and4_1 _11334_ (.A(net588),
    .B(net613),
    .C(net816),
    .D(net835),
    .X(_02129_));
 sky130_fd_sc_hd__nand2_4 _11335_ (.A(net602),
    .B(net827),
    .Y(_02130_));
 sky130_fd_sc_hd__a22oi_4 _11336_ (.A1(net613),
    .A2(net816),
    .B1(net835),
    .B2(net589),
    .Y(_02131_));
 sky130_fd_sc_hd__nor2_2 _11337_ (.A(_02129_),
    .B(_02131_),
    .Y(_02132_));
 sky130_fd_sc_hd__o21ba_4 _11338_ (.A1(_02130_),
    .A2(_02131_),
    .B1_N(_02129_),
    .X(_02133_));
 sky130_fd_sc_hd__nand2b_4 _11339_ (.A_N(_02133_),
    .B(_02128_),
    .Y(_02134_));
 sky130_fd_sc_hd__xnor2_4 _11340_ (.A(_02128_),
    .B(_02133_),
    .Y(_02135_));
 sky130_fd_sc_hd__and3_4 _11341_ (.A(_02125_),
    .B(_02126_),
    .C(_02135_),
    .X(_02136_));
 sky130_fd_sc_hd__o211ai_4 _11342_ (.A1(_02124_),
    .A2(_02136_),
    .B1(_02106_),
    .C1(_02107_),
    .Y(_02137_));
 sky130_fd_sc_hd__and2_1 _11343_ (.A(_02106_),
    .B(_02137_),
    .X(_02138_));
 sky130_fd_sc_hd__or2_1 _11344_ (.A(_02077_),
    .B(_02138_),
    .X(_02139_));
 sky130_fd_sc_hd__xor2_4 _11345_ (.A(_02089_),
    .B(_02090_),
    .X(_02140_));
 sky130_fd_sc_hd__a211o_2 _11346_ (.A1(_02106_),
    .A2(_02107_),
    .B1(_02124_),
    .C1(_02136_),
    .X(_02141_));
 sky130_fd_sc_hd__nand2_1 _11347_ (.A(_01698_),
    .B(_02045_),
    .Y(_02142_));
 sky130_fd_sc_hd__and2_2 _11348_ (.A(_02046_),
    .B(_02142_),
    .X(_02143_));
 sky130_fd_sc_hd__and3_2 _11349_ (.A(_02137_),
    .B(_02141_),
    .C(_02143_),
    .X(_02144_));
 sky130_fd_sc_hd__a21o_1 _11350_ (.A1(_02081_),
    .A2(_02082_),
    .B1(_02048_),
    .X(_02145_));
 sky130_fd_sc_hd__and3_1 _11351_ (.A(_02083_),
    .B(_02144_),
    .C(_02145_),
    .X(_02146_));
 sky130_fd_sc_hd__xnor2_2 _11352_ (.A(_02077_),
    .B(_02138_),
    .Y(_02147_));
 sky130_fd_sc_hd__a21oi_2 _11353_ (.A1(_02083_),
    .A2(_02145_),
    .B1(_02144_),
    .Y(_02148_));
 sky130_fd_sc_hd__or3_4 _11354_ (.A(_02146_),
    .B(_02147_),
    .C(_02148_),
    .X(_02149_));
 sky130_fd_sc_hd__nand2b_2 _11355_ (.A_N(_02146_),
    .B(_02149_),
    .Y(_02150_));
 sky130_fd_sc_hd__and2b_1 _11356_ (.A_N(_02140_),
    .B(_02150_),
    .X(_02151_));
 sky130_fd_sc_hd__xor2_2 _11357_ (.A(_02140_),
    .B(_02150_),
    .X(_02152_));
 sky130_fd_sc_hd__nor2_2 _11358_ (.A(_02139_),
    .B(_02152_),
    .Y(_02153_));
 sky130_fd_sc_hd__and2_2 _11359_ (.A(_02139_),
    .B(_02152_),
    .X(_02154_));
 sky130_fd_sc_hd__o21ai_2 _11360_ (.A1(_02146_),
    .A2(_02148_),
    .B1(_02147_),
    .Y(_02155_));
 sky130_fd_sc_hd__nand2_4 _11361_ (.A(_02149_),
    .B(_02155_),
    .Y(_02156_));
 sky130_fd_sc_hd__xnor2_4 _11362_ (.A(_02110_),
    .B(_02112_),
    .Y(_02157_));
 sky130_fd_sc_hd__nand2b_1 _11363_ (.A_N(_02034_),
    .B(_02157_),
    .Y(_02158_));
 sky130_fd_sc_hd__xnor2_1 _11364_ (.A(_02099_),
    .B(_02101_),
    .Y(_02159_));
 sky130_fd_sc_hd__or2_2 _11365_ (.A(_02158_),
    .B(_02159_),
    .X(_02160_));
 sky130_fd_sc_hd__a21oi_4 _11366_ (.A1(_02125_),
    .A2(_02126_),
    .B1(_02135_),
    .Y(_02161_));
 sky130_fd_sc_hd__or3_4 _11367_ (.A(_02136_),
    .B(_02160_),
    .C(_02161_),
    .X(_02162_));
 sky130_fd_sc_hd__o21ai_4 _11368_ (.A1(_02136_),
    .A2(_02161_),
    .B1(_02160_),
    .Y(_02163_));
 sky130_fd_sc_hd__xnor2_4 _11369_ (.A(_02120_),
    .B(_02122_),
    .Y(_02164_));
 sky130_fd_sc_hd__and4_1 _11370_ (.A(net515),
    .B(net523),
    .C(net907),
    .D(net916),
    .X(_02165_));
 sky130_fd_sc_hd__nand2_1 _11371_ (.A(net532),
    .B(net900),
    .Y(_02166_));
 sky130_fd_sc_hd__a22o_1 _11372_ (.A1(net523),
    .A2(net907),
    .B1(net916),
    .B2(net515),
    .X(_02167_));
 sky130_fd_sc_hd__and2b_1 _11373_ (.A_N(_02165_),
    .B(_02167_),
    .X(_02168_));
 sky130_fd_sc_hd__a31o_2 _11374_ (.A1(net532),
    .A2(net900),
    .A3(_02167_),
    .B1(_02165_),
    .X(_02169_));
 sky130_fd_sc_hd__a22o_2 _11375_ (.A1(net578),
    .A2(net856),
    .B1(_02117_),
    .B2(_02118_),
    .X(_02170_));
 sky130_fd_sc_hd__nand3_4 _11376_ (.A(_02119_),
    .B(_02169_),
    .C(_02170_),
    .Y(_02171_));
 sky130_fd_sc_hd__and4_1 _11377_ (.A(net545),
    .B(net561),
    .C(net877),
    .D(net887),
    .X(_02172_));
 sky130_fd_sc_hd__nand2_1 _11378_ (.A(net578),
    .B(net866),
    .Y(_02173_));
 sky130_fd_sc_hd__a22oi_4 _11379_ (.A1(net561),
    .A2(net877),
    .B1(net887),
    .B2(net545),
    .Y(_02174_));
 sky130_fd_sc_hd__or3_2 _11380_ (.A(_02172_),
    .B(_02173_),
    .C(_02174_),
    .X(_02175_));
 sky130_fd_sc_hd__nand2b_2 _11381_ (.A_N(_02172_),
    .B(_02175_),
    .Y(_02176_));
 sky130_fd_sc_hd__a21o_1 _11382_ (.A1(_02119_),
    .A2(_02170_),
    .B1(_02169_),
    .X(_02177_));
 sky130_fd_sc_hd__nand3_4 _11383_ (.A(_02171_),
    .B(_02176_),
    .C(_02177_),
    .Y(_02178_));
 sky130_fd_sc_hd__a21oi_4 _11384_ (.A1(_02171_),
    .A2(_02178_),
    .B1(_02164_),
    .Y(_02179_));
 sky130_fd_sc_hd__a21o_1 _11385_ (.A1(_02171_),
    .A2(_02178_),
    .B1(_02164_),
    .X(_02180_));
 sky130_fd_sc_hd__xnor2_4 _11386_ (.A(_02130_),
    .B(_02132_),
    .Y(_02181_));
 sky130_fd_sc_hd__and3_2 _11387_ (.A(net590),
    .B(net846),
    .C(_02072_),
    .X(_02182_));
 sky130_fd_sc_hd__nand2_2 _11388_ (.A(net604),
    .B(net835),
    .Y(_02183_));
 sky130_fd_sc_hd__and2_1 _11389_ (.A(net590),
    .B(net846),
    .X(_02184_));
 sky130_fd_sc_hd__o21ba_2 _11390_ (.A1(_02072_),
    .A2(_02184_),
    .B1_N(_02182_),
    .X(_02185_));
 sky130_fd_sc_hd__and3_1 _11391_ (.A(net602),
    .B(net835),
    .C(_02185_),
    .X(_02186_));
 sky130_fd_sc_hd__o21ai_4 _11392_ (.A1(_02182_),
    .A2(_02186_),
    .B1(_02181_),
    .Y(_02187_));
 sky130_fd_sc_hd__or3_1 _11393_ (.A(_02181_),
    .B(_02182_),
    .C(_02186_),
    .X(_02188_));
 sky130_fd_sc_hd__and2_2 _11394_ (.A(_02187_),
    .B(_02188_),
    .X(_02189_));
 sky130_fd_sc_hd__nand3_2 _11395_ (.A(_02164_),
    .B(_02171_),
    .C(_02178_),
    .Y(_02190_));
 sky130_fd_sc_hd__and3_4 _11396_ (.A(_02180_),
    .B(_02189_),
    .C(_02190_),
    .X(_02191_));
 sky130_fd_sc_hd__o211ai_4 _11397_ (.A1(_02179_),
    .A2(_02191_),
    .B1(_02162_),
    .C1(_02163_),
    .Y(_02192_));
 sky130_fd_sc_hd__a211o_2 _11398_ (.A1(_02162_),
    .A2(_02163_),
    .B1(_02179_),
    .C1(_02191_),
    .X(_02193_));
 sky130_fd_sc_hd__xnor2_4 _11399_ (.A(_02102_),
    .B(_02103_),
    .Y(_02194_));
 sky130_fd_sc_hd__and3_2 _11400_ (.A(_02192_),
    .B(_02193_),
    .C(_02194_),
    .X(_02195_));
 sky130_fd_sc_hd__a21oi_4 _11401_ (.A1(_02137_),
    .A2(_02141_),
    .B1(_02143_),
    .Y(_02196_));
 sky130_fd_sc_hd__nor3b_4 _11402_ (.A(_02144_),
    .B(_02196_),
    .C_N(_02195_),
    .Y(_02197_));
 sky130_fd_sc_hd__and2_2 _11403_ (.A(_02162_),
    .B(_02192_),
    .X(_02198_));
 sky130_fd_sc_hd__or2_1 _11404_ (.A(_02134_),
    .B(_02198_),
    .X(_02199_));
 sky130_fd_sc_hd__inv_2 _11405_ (.A(_02199_),
    .Y(_02200_));
 sky130_fd_sc_hd__xnor2_4 _11406_ (.A(_02134_),
    .B(_02198_),
    .Y(_02201_));
 sky130_fd_sc_hd__o21ba_2 _11407_ (.A1(_02144_),
    .A2(_02196_),
    .B1_N(_02195_),
    .X(_02202_));
 sky130_fd_sc_hd__or3_4 _11408_ (.A(_02197_),
    .B(_02201_),
    .C(_02202_),
    .X(_02203_));
 sky130_fd_sc_hd__and2b_2 _11409_ (.A_N(_02197_),
    .B(_02203_),
    .X(_02204_));
 sky130_fd_sc_hd__nor2_1 _11410_ (.A(_02156_),
    .B(_02204_),
    .Y(_02205_));
 sky130_fd_sc_hd__xor2_4 _11411_ (.A(_02156_),
    .B(_02204_),
    .X(_02206_));
 sky130_fd_sc_hd__a21oi_2 _11412_ (.A1(_02200_),
    .A2(_02206_),
    .B1(_02205_),
    .Y(_02207_));
 sky130_fd_sc_hd__nor3_4 _11413_ (.A(_02153_),
    .B(_02154_),
    .C(_02207_),
    .Y(_02208_));
 sky130_fd_sc_hd__o21ai_2 _11414_ (.A1(_02092_),
    .A2(_02093_),
    .B1(_02087_),
    .Y(_02209_));
 sky130_fd_sc_hd__nand2_4 _11415_ (.A(_02094_),
    .B(_02209_),
    .Y(_02210_));
 sky130_fd_sc_hd__or2_4 _11416_ (.A(_02151_),
    .B(_02153_),
    .X(_02211_));
 sky130_fd_sc_hd__and2b_2 _11417_ (.A_N(_02210_),
    .B(_02211_),
    .X(_02212_));
 sky130_fd_sc_hd__xnor2_4 _11418_ (.A(_02210_),
    .B(_02211_),
    .Y(_02213_));
 sky130_fd_sc_hd__xnor2_4 _11419_ (.A(_02200_),
    .B(_02206_),
    .Y(_02214_));
 sky130_fd_sc_hd__o21ai_4 _11420_ (.A1(_02197_),
    .A2(_02202_),
    .B1(_02201_),
    .Y(_02215_));
 sky130_fd_sc_hd__a21oi_4 _11421_ (.A1(_02180_),
    .A2(_02190_),
    .B1(_02189_),
    .Y(_02216_));
 sky130_fd_sc_hd__a21o_1 _11422_ (.A1(_02171_),
    .A2(_02177_),
    .B1(_02176_),
    .X(_02217_));
 sky130_fd_sc_hd__and4_2 _11423_ (.A(net522),
    .B(net532),
    .C(net907),
    .D(net916),
    .X(_02218_));
 sky130_fd_sc_hd__inv_2 _11424_ (.A(_02218_),
    .Y(_02219_));
 sky130_fd_sc_hd__o21ai_2 _11425_ (.A1(_02172_),
    .A2(_02174_),
    .B1(_02173_),
    .Y(_02220_));
 sky130_fd_sc_hd__nand3_2 _11426_ (.A(_02175_),
    .B(_02218_),
    .C(_02220_),
    .Y(_02221_));
 sky130_fd_sc_hd__and4_2 _11427_ (.A(net546),
    .B(net561),
    .C(net887),
    .D(net897),
    .X(_02222_));
 sky130_fd_sc_hd__nand2_2 _11428_ (.A(net578),
    .B(net876),
    .Y(_02223_));
 sky130_fd_sc_hd__a22oi_4 _11429_ (.A1(net561),
    .A2(net887),
    .B1(net897),
    .B2(net546),
    .Y(_02224_));
 sky130_fd_sc_hd__or3_4 _11430_ (.A(_02222_),
    .B(_02223_),
    .C(_02224_),
    .X(_02225_));
 sky130_fd_sc_hd__nand2b_2 _11431_ (.A_N(_02222_),
    .B(_02225_),
    .Y(_02226_));
 sky130_fd_sc_hd__a21o_1 _11432_ (.A1(_02175_),
    .A2(_02220_),
    .B1(_02218_),
    .X(_02227_));
 sky130_fd_sc_hd__nand3_2 _11433_ (.A(_02221_),
    .B(_02226_),
    .C(_02227_),
    .Y(_02228_));
 sky130_fd_sc_hd__a21bo_2 _11434_ (.A1(_02226_),
    .A2(_02227_),
    .B1_N(_02221_),
    .X(_02229_));
 sky130_fd_sc_hd__nand3_4 _11435_ (.A(_02178_),
    .B(_02217_),
    .C(_02229_),
    .Y(_02230_));
 sky130_fd_sc_hd__xnor2_4 _11436_ (.A(_02183_),
    .B(_02185_),
    .Y(_02231_));
 sky130_fd_sc_hd__and4_2 _11437_ (.A(net591),
    .B(net614),
    .C(net836),
    .D(net856),
    .X(_02232_));
 sky130_fd_sc_hd__a22oi_2 _11438_ (.A1(net614),
    .A2(net836),
    .B1(net857),
    .B2(net591),
    .Y(_02233_));
 sky130_fd_sc_hd__and4bb_2 _11439_ (.A_N(_02232_),
    .B_N(_02233_),
    .C(net603),
    .D(net847),
    .X(_02234_));
 sky130_fd_sc_hd__nor2_4 _11440_ (.A(_02232_),
    .B(_02234_),
    .Y(_02235_));
 sky130_fd_sc_hd__nand2b_1 _11441_ (.A_N(_02235_),
    .B(_02231_),
    .Y(_02236_));
 sky130_fd_sc_hd__xnor2_4 _11442_ (.A(_02231_),
    .B(_02235_),
    .Y(_02237_));
 sky130_fd_sc_hd__a21o_1 _11443_ (.A1(_02178_),
    .A2(_02217_),
    .B1(_02229_),
    .X(_02238_));
 sky130_fd_sc_hd__nand3_4 _11444_ (.A(_02230_),
    .B(_02237_),
    .C(_02238_),
    .Y(_02239_));
 sky130_fd_sc_hd__a211o_2 _11445_ (.A1(_02230_),
    .A2(_02239_),
    .B1(_02191_),
    .C1(_02216_),
    .X(_02240_));
 sky130_fd_sc_hd__o211ai_4 _11446_ (.A1(_02191_),
    .A2(_02216_),
    .B1(_02230_),
    .C1(_02239_),
    .Y(_02241_));
 sky130_fd_sc_hd__nand2_1 _11447_ (.A(_02158_),
    .B(_02159_),
    .Y(_02242_));
 sky130_fd_sc_hd__and2_2 _11448_ (.A(_02160_),
    .B(_02242_),
    .X(_02243_));
 sky130_fd_sc_hd__and3_2 _11449_ (.A(_02240_),
    .B(_02241_),
    .C(_02243_),
    .X(_02244_));
 sky130_fd_sc_hd__a21oi_4 _11450_ (.A1(_02192_),
    .A2(_02193_),
    .B1(_02194_),
    .Y(_02245_));
 sky130_fd_sc_hd__nor3b_4 _11451_ (.A(_02195_),
    .B(_02245_),
    .C_N(_02244_),
    .Y(_02246_));
 sky130_fd_sc_hd__or2_4 _11452_ (.A(_02187_),
    .B(_02240_),
    .X(_02247_));
 sky130_fd_sc_hd__nand2_1 _11453_ (.A(_02187_),
    .B(_02240_),
    .Y(_02248_));
 sky130_fd_sc_hd__nand2_4 _11454_ (.A(_02247_),
    .B(_02248_),
    .Y(_02249_));
 sky130_fd_sc_hd__o21ba_4 _11455_ (.A1(_02195_),
    .A2(_02245_),
    .B1_N(_02244_),
    .X(_02250_));
 sky130_fd_sc_hd__or3_4 _11456_ (.A(_02246_),
    .B(_02249_),
    .C(_02250_),
    .X(_02251_));
 sky130_fd_sc_hd__o21bai_4 _11457_ (.A1(_02249_),
    .A2(_02250_),
    .B1_N(_02246_),
    .Y(_02252_));
 sky130_fd_sc_hd__and3_2 _11458_ (.A(_02203_),
    .B(_02215_),
    .C(_02252_),
    .X(_02253_));
 sky130_fd_sc_hd__a21oi_4 _11459_ (.A1(_02203_),
    .A2(_02215_),
    .B1(_02252_),
    .Y(_02254_));
 sky130_fd_sc_hd__or3_4 _11460_ (.A(_02247_),
    .B(_02253_),
    .C(_02254_),
    .X(_02255_));
 sky130_fd_sc_hd__and2b_2 _11461_ (.A_N(_02253_),
    .B(_02255_),
    .X(_02256_));
 sky130_fd_sc_hd__or2_4 _11462_ (.A(_02214_),
    .B(_02256_),
    .X(_02257_));
 sky130_fd_sc_hd__o21a_1 _11463_ (.A1(_02153_),
    .A2(_02154_),
    .B1(_02207_),
    .X(_02258_));
 sky130_fd_sc_hd__or2_4 _11464_ (.A(_02208_),
    .B(_02258_),
    .X(_02259_));
 sky130_fd_sc_hd__xor2_4 _11465_ (.A(_02257_),
    .B(_02259_),
    .X(_02260_));
 sky130_fd_sc_hd__a21o_1 _11466_ (.A1(_02230_),
    .A2(_02238_),
    .B1(_02237_),
    .X(_02261_));
 sky130_fd_sc_hd__and4_1 _11467_ (.A(net545),
    .B(net560),
    .C(net897),
    .D(net905),
    .X(_02262_));
 sky130_fd_sc_hd__nand4_1 _11468_ (.A(net545),
    .B(net560),
    .C(net897),
    .D(net905),
    .Y(_02263_));
 sky130_fd_sc_hd__and2_2 _11469_ (.A(net578),
    .B(net887),
    .X(_02264_));
 sky130_fd_sc_hd__nand2_1 _11470_ (.A(net578),
    .B(net887),
    .Y(_02265_));
 sky130_fd_sc_hd__a22o_1 _11471_ (.A1(net560),
    .A2(net898),
    .B1(net905),
    .B2(net545),
    .X(_02266_));
 sky130_fd_sc_hd__or3b_4 _11472_ (.A(_02262_),
    .B(_02265_),
    .C_N(_02266_),
    .X(_02267_));
 sky130_fd_sc_hd__a21o_2 _11473_ (.A1(_02264_),
    .A2(_02266_),
    .B1(_02262_),
    .X(_02268_));
 sky130_fd_sc_hd__o21ai_4 _11474_ (.A1(_02222_),
    .A2(_02224_),
    .B1(_02223_),
    .Y(_02269_));
 sky130_fd_sc_hd__and3_4 _11475_ (.A(_02225_),
    .B(_02268_),
    .C(_02269_),
    .X(_02270_));
 sky130_fd_sc_hd__a21o_2 _11476_ (.A1(_02221_),
    .A2(_02227_),
    .B1(_02226_),
    .X(_02271_));
 sky130_fd_sc_hd__and3_4 _11477_ (.A(_02228_),
    .B(_02270_),
    .C(_02271_),
    .X(_02272_));
 sky130_fd_sc_hd__o2bb2a_1 _11478_ (.A1_N(net604),
    .A2_N(net846),
    .B1(_02232_),
    .B2(_02233_),
    .X(_02273_));
 sky130_fd_sc_hd__nor2_1 _11479_ (.A(_02234_),
    .B(_02273_),
    .Y(_02274_));
 sky130_fd_sc_hd__and4_2 _11480_ (.A(net591),
    .B(net614),
    .C(net848),
    .D(net867),
    .X(_02275_));
 sky130_fd_sc_hd__a22oi_2 _11481_ (.A1(net614),
    .A2(net848),
    .B1(net867),
    .B2(net590),
    .Y(_02276_));
 sky130_fd_sc_hd__and4bb_2 _11482_ (.A_N(_02275_),
    .B_N(_02276_),
    .C(net603),
    .D(net858),
    .X(_02277_));
 sky130_fd_sc_hd__o21ai_2 _11483_ (.A1(_02275_),
    .A2(_02277_),
    .B1(_02274_),
    .Y(_02278_));
 sky130_fd_sc_hd__or3_1 _11484_ (.A(_02274_),
    .B(_02275_),
    .C(_02277_),
    .X(_02279_));
 sky130_fd_sc_hd__and2_1 _11485_ (.A(_02278_),
    .B(_02279_),
    .X(_02280_));
 sky130_fd_sc_hd__a21oi_4 _11486_ (.A1(_02228_),
    .A2(_02271_),
    .B1(_02270_),
    .Y(_02281_));
 sky130_fd_sc_hd__nor3b_4 _11487_ (.A(_02272_),
    .B(_02281_),
    .C_N(_02280_),
    .Y(_02282_));
 sky130_fd_sc_hd__o211ai_4 _11488_ (.A1(_02272_),
    .A2(_02282_),
    .B1(_02239_),
    .C1(_02261_),
    .Y(_02283_));
 sky130_fd_sc_hd__or2_4 _11489_ (.A(_02236_),
    .B(_02283_),
    .X(_02284_));
 sky130_fd_sc_hd__o21ai_4 _11490_ (.A1(_02246_),
    .A2(_02250_),
    .B1(_02249_),
    .Y(_02285_));
 sky130_fd_sc_hd__a211o_2 _11491_ (.A1(_02239_),
    .A2(_02261_),
    .B1(_02272_),
    .C1(_02282_),
    .X(_02286_));
 sky130_fd_sc_hd__xnor2_4 _11492_ (.A(_02034_),
    .B(_02157_),
    .Y(_02287_));
 sky130_fd_sc_hd__and3_2 _11493_ (.A(_02283_),
    .B(_02286_),
    .C(_02287_),
    .X(_02288_));
 sky130_fd_sc_hd__a21oi_4 _11494_ (.A1(_02240_),
    .A2(_02241_),
    .B1(_02243_),
    .Y(_02289_));
 sky130_fd_sc_hd__nor3b_4 _11495_ (.A(_02244_),
    .B(_02289_),
    .C_N(_02288_),
    .Y(_02290_));
 sky130_fd_sc_hd__nand2_1 _11496_ (.A(_02236_),
    .B(_02283_),
    .Y(_02291_));
 sky130_fd_sc_hd__nand2_2 _11497_ (.A(_02284_),
    .B(_02291_),
    .Y(_02292_));
 sky130_fd_sc_hd__o21ba_2 _11498_ (.A1(_02244_),
    .A2(_02289_),
    .B1_N(_02288_),
    .X(_02293_));
 sky130_fd_sc_hd__nor3_4 _11499_ (.A(_02290_),
    .B(_02292_),
    .C(_02293_),
    .Y(_02294_));
 sky130_fd_sc_hd__o211a_4 _11500_ (.A1(_02290_),
    .A2(_02294_),
    .B1(_02251_),
    .C1(_02285_),
    .X(_02295_));
 sky130_fd_sc_hd__a211oi_4 _11501_ (.A1(_02251_),
    .A2(_02285_),
    .B1(_02290_),
    .C1(_02294_),
    .Y(_02296_));
 sky130_fd_sc_hd__nor3_4 _11502_ (.A(_02284_),
    .B(_02295_),
    .C(_02296_),
    .Y(_02297_));
 sky130_fd_sc_hd__o21a_1 _11503_ (.A1(_02295_),
    .A2(_02296_),
    .B1(_02284_),
    .X(_02298_));
 sky130_fd_sc_hd__o21a_2 _11504_ (.A1(_02290_),
    .A2(_02293_),
    .B1(_02292_),
    .X(_02299_));
 sky130_fd_sc_hd__o21ba_2 _11505_ (.A1(_02272_),
    .A2(_02281_),
    .B1_N(_02280_),
    .X(_02300_));
 sky130_fd_sc_hd__and4_1 _11506_ (.A(net545),
    .B(net560),
    .C(net907),
    .D(net914),
    .X(_02301_));
 sky130_fd_sc_hd__a22oi_1 _11507_ (.A1(net560),
    .A2(net907),
    .B1(net914),
    .B2(net545),
    .Y(_02302_));
 sky130_fd_sc_hd__a22o_1 _11508_ (.A1(net560),
    .A2(net907),
    .B1(net914),
    .B2(net545),
    .X(_02303_));
 sky130_fd_sc_hd__and4b_1 _11509_ (.A_N(_02301_),
    .B(_02303_),
    .C(net578),
    .D(net898),
    .X(_02304_));
 sky130_fd_sc_hd__a31o_2 _11510_ (.A1(net578),
    .A2(net898),
    .A3(_02303_),
    .B1(_02301_),
    .X(_02305_));
 sky130_fd_sc_hd__a21o_1 _11511_ (.A1(_02263_),
    .A2(_02266_),
    .B1(_02264_),
    .X(_02306_));
 sky130_fd_sc_hd__nand3_4 _11512_ (.A(_02267_),
    .B(_02305_),
    .C(_02306_),
    .Y(_02307_));
 sky130_fd_sc_hd__a21oi_4 _11513_ (.A1(_02225_),
    .A2(_02269_),
    .B1(_02268_),
    .Y(_02308_));
 sky130_fd_sc_hd__or3_4 _11514_ (.A(_02270_),
    .B(_02307_),
    .C(_02308_),
    .X(_02309_));
 sky130_fd_sc_hd__o2bb2a_1 _11515_ (.A1_N(net603),
    .A2_N(net858),
    .B1(_02275_),
    .B2(_02276_),
    .X(_02310_));
 sky130_fd_sc_hd__nor2_2 _11516_ (.A(_02277_),
    .B(_02310_),
    .Y(_02311_));
 sky130_fd_sc_hd__nand2_4 _11517_ (.A(net614),
    .B(net876),
    .Y(_02312_));
 sky130_fd_sc_hd__and4_2 _11518_ (.A(net590),
    .B(net612),
    .C(net857),
    .D(net876),
    .X(_02313_));
 sky130_fd_sc_hd__a22oi_2 _11519_ (.A1(net613),
    .A2(net857),
    .B1(net877),
    .B2(net590),
    .Y(_02314_));
 sky130_fd_sc_hd__and4bb_2 _11520_ (.A_N(_02313_),
    .B_N(_02314_),
    .C(net602),
    .D(net866),
    .X(_02315_));
 sky130_fd_sc_hd__nor2_4 _11521_ (.A(_02313_),
    .B(_02315_),
    .Y(_02316_));
 sky130_fd_sc_hd__or3_2 _11522_ (.A(_02277_),
    .B(_02310_),
    .C(_02316_),
    .X(_02317_));
 sky130_fd_sc_hd__xnor2_4 _11523_ (.A(_02311_),
    .B(_02316_),
    .Y(_02318_));
 sky130_fd_sc_hd__o21ai_4 _11524_ (.A1(_02270_),
    .A2(_02308_),
    .B1(_02307_),
    .Y(_02319_));
 sky130_fd_sc_hd__nand3_4 _11525_ (.A(_02309_),
    .B(_02318_),
    .C(_02319_),
    .Y(_02320_));
 sky130_fd_sc_hd__nand2_1 _11526_ (.A(_02309_),
    .B(_02320_),
    .Y(_02321_));
 sky130_fd_sc_hd__or3b_4 _11527_ (.A(_02282_),
    .B(_02300_),
    .C_N(_02321_),
    .X(_02322_));
 sky130_fd_sc_hd__o21bai_4 _11528_ (.A1(_02282_),
    .A2(_02300_),
    .B1_N(_02321_),
    .Y(_02323_));
 sky130_fd_sc_hd__xnor2_2 _11529_ (.A(_02166_),
    .B(_02168_),
    .Y(_02324_));
 sky130_fd_sc_hd__and3_2 _11530_ (.A(_02322_),
    .B(_02323_),
    .C(_02324_),
    .X(_02325_));
 sky130_fd_sc_hd__a21oi_4 _11531_ (.A1(_02283_),
    .A2(_02286_),
    .B1(_02287_),
    .Y(_02326_));
 sky130_fd_sc_hd__nor3b_4 _11532_ (.A(_02288_),
    .B(_02326_),
    .C_N(_02325_),
    .Y(_02327_));
 sky130_fd_sc_hd__or2_4 _11533_ (.A(_02278_),
    .B(_02322_),
    .X(_02328_));
 sky130_fd_sc_hd__nand2_1 _11534_ (.A(_02278_),
    .B(_02322_),
    .Y(_02329_));
 sky130_fd_sc_hd__nand2_2 _11535_ (.A(_02328_),
    .B(_02329_),
    .Y(_02330_));
 sky130_fd_sc_hd__o21ba_2 _11536_ (.A1(_02288_),
    .A2(_02326_),
    .B1_N(_02325_),
    .X(_02331_));
 sky130_fd_sc_hd__nor3_4 _11537_ (.A(_02327_),
    .B(_02330_),
    .C(_02331_),
    .Y(_02332_));
 sky130_fd_sc_hd__or2_1 _11538_ (.A(_02327_),
    .B(_02332_),
    .X(_02333_));
 sky130_fd_sc_hd__nor3b_4 _11539_ (.A(_02294_),
    .B(_02299_),
    .C_N(_02333_),
    .Y(_02334_));
 sky130_fd_sc_hd__o21ba_2 _11540_ (.A1(_02294_),
    .A2(_02299_),
    .B1_N(_02333_),
    .X(_02335_));
 sky130_fd_sc_hd__nor3_4 _11541_ (.A(_02328_),
    .B(_02334_),
    .C(_02335_),
    .Y(_02336_));
 sky130_fd_sc_hd__or2_1 _11542_ (.A(_02334_),
    .B(_02336_),
    .X(_02337_));
 sky130_fd_sc_hd__or3b_2 _11543_ (.A(_02297_),
    .B(_02298_),
    .C_N(_02337_),
    .X(_02338_));
 sky130_fd_sc_hd__o21ai_4 _11544_ (.A1(_02253_),
    .A2(_02254_),
    .B1(_02247_),
    .Y(_02339_));
 sky130_fd_sc_hd__o211ai_4 _11545_ (.A1(_02295_),
    .A2(_02297_),
    .B1(_02339_),
    .C1(_02255_),
    .Y(_02340_));
 sky130_fd_sc_hd__a211o_1 _11546_ (.A1(_02255_),
    .A2(_02339_),
    .B1(_02297_),
    .C1(_02295_),
    .X(_02341_));
 sky130_fd_sc_hd__nand3b_2 _11547_ (.A_N(_02338_),
    .B(_02340_),
    .C(_02341_),
    .Y(_02342_));
 sky130_fd_sc_hd__a21bo_1 _11548_ (.A1(_02340_),
    .A2(_02341_),
    .B1_N(_02338_),
    .X(_02343_));
 sky130_fd_sc_hd__and2_1 _11549_ (.A(_02342_),
    .B(_02343_),
    .X(_02344_));
 sky130_fd_sc_hd__o21a_2 _11550_ (.A1(_02334_),
    .A2(_02335_),
    .B1(_02328_),
    .X(_02345_));
 sky130_fd_sc_hd__o21a_2 _11551_ (.A1(_02327_),
    .A2(_02331_),
    .B1(_02330_),
    .X(_02346_));
 sky130_fd_sc_hd__a21o_1 _11552_ (.A1(_02309_),
    .A2(_02319_),
    .B1(_02318_),
    .X(_02347_));
 sky130_fd_sc_hd__and4_1 _11553_ (.A(net562),
    .B(net579),
    .C(net907),
    .D(net917),
    .X(_02348_));
 sky130_fd_sc_hd__o22a_1 _11554_ (.A1(net304),
    .A2(_03280_),
    .B1(_02301_),
    .B2(_02302_),
    .X(_02349_));
 sky130_fd_sc_hd__nor3b_2 _11555_ (.A(_02304_),
    .B(_02349_),
    .C_N(_02348_),
    .Y(_02350_));
 sky130_fd_sc_hd__a21o_1 _11556_ (.A1(_02267_),
    .A2(_02306_),
    .B1(_02305_),
    .X(_02351_));
 sky130_fd_sc_hd__and3_2 _11557_ (.A(_02307_),
    .B(_02350_),
    .C(_02351_),
    .X(_02352_));
 sky130_fd_sc_hd__nand3_1 _11558_ (.A(_02307_),
    .B(_02350_),
    .C(_02351_),
    .Y(_02353_));
 sky130_fd_sc_hd__o2bb2a_1 _11559_ (.A1_N(net602),
    .A2_N(net865),
    .B1(_02313_),
    .B2(_02314_),
    .X(_02354_));
 sky130_fd_sc_hd__nor2_1 _11560_ (.A(_02315_),
    .B(_02354_),
    .Y(_02355_));
 sky130_fd_sc_hd__and4_1 _11561_ (.A(net590),
    .B(net612),
    .C(net865),
    .D(net887),
    .X(_02356_));
 sky130_fd_sc_hd__a22oi_2 _11562_ (.A1(net612),
    .A2(net865),
    .B1(net887),
    .B2(net590),
    .Y(_02357_));
 sky130_fd_sc_hd__and4bb_2 _11563_ (.A_N(_02356_),
    .B_N(_02357_),
    .C(net602),
    .D(net876),
    .X(_02358_));
 sky130_fd_sc_hd__nor2_1 _11564_ (.A(_02356_),
    .B(_02358_),
    .Y(_02359_));
 sky130_fd_sc_hd__or3_2 _11565_ (.A(_02315_),
    .B(_02354_),
    .C(_02359_),
    .X(_02360_));
 sky130_fd_sc_hd__xnor2_1 _11566_ (.A(_02355_),
    .B(_02359_),
    .Y(_02361_));
 sky130_fd_sc_hd__a21o_1 _11567_ (.A1(_02307_),
    .A2(_02351_),
    .B1(_02350_),
    .X(_02362_));
 sky130_fd_sc_hd__and3_2 _11568_ (.A(_02353_),
    .B(_02361_),
    .C(_02362_),
    .X(_02363_));
 sky130_fd_sc_hd__o211ai_4 _11569_ (.A1(_02352_),
    .A2(_02363_),
    .B1(_02320_),
    .C1(_02347_),
    .Y(_02364_));
 sky130_fd_sc_hd__a211o_2 _11570_ (.A1(_02320_),
    .A2(_02347_),
    .B1(_02352_),
    .C1(_02363_),
    .X(_02365_));
 sky130_fd_sc_hd__a22o_2 _11571_ (.A1(net532),
    .A2(net907),
    .B1(net917),
    .B2(net522),
    .X(_02366_));
 sky130_fd_sc_hd__nand4_4 _11572_ (.A(_02219_),
    .B(_02364_),
    .C(_02365_),
    .D(_02366_),
    .Y(_02367_));
 sky130_fd_sc_hd__a21oi_4 _11573_ (.A1(_02322_),
    .A2(_02323_),
    .B1(_02324_),
    .Y(_02368_));
 sky130_fd_sc_hd__or3_4 _11574_ (.A(_02325_),
    .B(_02367_),
    .C(_02368_),
    .X(_02369_));
 sky130_fd_sc_hd__nor2_4 _11575_ (.A(_02317_),
    .B(_02364_),
    .Y(_02370_));
 sky130_fd_sc_hd__and2_1 _11576_ (.A(_02317_),
    .B(_02364_),
    .X(_02371_));
 sky130_fd_sc_hd__nor2_2 _11577_ (.A(_02370_),
    .B(_02371_),
    .Y(_02372_));
 sky130_fd_sc_hd__o21ai_4 _11578_ (.A1(_02325_),
    .A2(_02368_),
    .B1(_02367_),
    .Y(_02373_));
 sky130_fd_sc_hd__nand3_4 _11579_ (.A(_02369_),
    .B(_02372_),
    .C(_02373_),
    .Y(_02374_));
 sky130_fd_sc_hd__a211o_2 _11580_ (.A1(_02369_),
    .A2(_02374_),
    .B1(_02332_),
    .C1(_02346_),
    .X(_02375_));
 sky130_fd_sc_hd__o211ai_4 _11581_ (.A1(_02332_),
    .A2(_02346_),
    .B1(_02369_),
    .C1(_02374_),
    .Y(_02376_));
 sky130_fd_sc_hd__nand3_4 _11582_ (.A(_02370_),
    .B(_02375_),
    .C(_02376_),
    .Y(_02377_));
 sky130_fd_sc_hd__nand2_1 _11583_ (.A(_02375_),
    .B(_02377_),
    .Y(_02378_));
 sky130_fd_sc_hd__nor3b_4 _11584_ (.A(_02336_),
    .B(_02345_),
    .C_N(_02378_),
    .Y(_02379_));
 sky130_fd_sc_hd__o21bai_1 _11585_ (.A1(_02297_),
    .A2(_02298_),
    .B1_N(_02337_),
    .Y(_02380_));
 sky130_fd_sc_hd__nand3_1 _11586_ (.A(_02338_),
    .B(_02379_),
    .C(_02380_),
    .Y(_02381_));
 sky130_fd_sc_hd__a21o_1 _11587_ (.A1(_02375_),
    .A2(_02376_),
    .B1(_02370_),
    .X(_02382_));
 sky130_fd_sc_hd__a21o_1 _11588_ (.A1(_02369_),
    .A2(_02373_),
    .B1(_02372_),
    .X(_02383_));
 sky130_fd_sc_hd__o2bb2a_1 _11589_ (.A1_N(net602),
    .A2_N(net876),
    .B1(_02356_),
    .B2(_02357_),
    .X(_02384_));
 sky130_fd_sc_hd__nor2_4 _11590_ (.A(_02358_),
    .B(_02384_),
    .Y(_02385_));
 sky130_fd_sc_hd__and2_4 _11591_ (.A(net590),
    .B(net898),
    .X(_02386_));
 sky130_fd_sc_hd__nand2_2 _11592_ (.A(net590),
    .B(net899),
    .Y(_02387_));
 sky130_fd_sc_hd__nor2_1 _11593_ (.A(_02312_),
    .B(_02387_),
    .Y(_02388_));
 sky130_fd_sc_hd__nand2_2 _11594_ (.A(net603),
    .B(net889),
    .Y(_02389_));
 sky130_fd_sc_hd__xnor2_4 _11595_ (.A(_02312_),
    .B(_02386_),
    .Y(_02390_));
 sky130_fd_sc_hd__a31o_4 _11596_ (.A1(net603),
    .A2(net889),
    .A3(_02390_),
    .B1(_02388_),
    .X(_02391_));
 sky130_fd_sc_hd__and2_4 _11597_ (.A(_02385_),
    .B(_02391_),
    .X(_02392_));
 sky130_fd_sc_hd__xor2_4 _11598_ (.A(_02385_),
    .B(_02391_),
    .X(_02393_));
 sky130_fd_sc_hd__o21bai_1 _11599_ (.A1(_02304_),
    .A2(_02349_),
    .B1_N(_02348_),
    .Y(_02394_));
 sky130_fd_sc_hd__and2b_1 _11600_ (.A_N(_02350_),
    .B(_02394_),
    .X(_02395_));
 sky130_fd_sc_hd__nand2_1 _11601_ (.A(_02393_),
    .B(_02395_),
    .Y(_02396_));
 sky130_fd_sc_hd__a21oi_1 _11602_ (.A1(_02353_),
    .A2(_02362_),
    .B1(_02361_),
    .Y(_02397_));
 sky130_fd_sc_hd__or3_2 _11603_ (.A(_02363_),
    .B(_02396_),
    .C(_02397_),
    .X(_02398_));
 sky130_fd_sc_hd__o21ai_1 _11604_ (.A1(_02363_),
    .A2(_02397_),
    .B1(_02396_),
    .Y(_02399_));
 sky130_fd_sc_hd__and4_1 _11605_ (.A(net533),
    .B(net917),
    .C(_02398_),
    .D(_02399_),
    .X(_02400_));
 sky130_fd_sc_hd__a22o_1 _11606_ (.A1(_02364_),
    .A2(_02365_),
    .B1(_02366_),
    .B2(_02219_),
    .X(_02401_));
 sky130_fd_sc_hd__nand3_1 _11607_ (.A(_02367_),
    .B(_02400_),
    .C(_02401_),
    .Y(_02402_));
 sky130_fd_sc_hd__a21o_1 _11608_ (.A1(_02367_),
    .A2(_02401_),
    .B1(_02400_),
    .X(_02403_));
 sky130_fd_sc_hd__or2_4 _11609_ (.A(_02360_),
    .B(_02398_),
    .X(_02404_));
 sky130_fd_sc_hd__nand2_1 _11610_ (.A(_02360_),
    .B(_02398_),
    .Y(_02405_));
 sky130_fd_sc_hd__and2_1 _11611_ (.A(_02404_),
    .B(_02405_),
    .X(_02406_));
 sky130_fd_sc_hd__nand3_1 _11612_ (.A(_02402_),
    .B(_02403_),
    .C(_02406_),
    .Y(_02407_));
 sky130_fd_sc_hd__nand2_1 _11613_ (.A(_02402_),
    .B(_02407_),
    .Y(_02408_));
 sky130_fd_sc_hd__and3_4 _11614_ (.A(_02374_),
    .B(_02383_),
    .C(_02408_),
    .X(_02409_));
 sky130_fd_sc_hd__a21oi_2 _11615_ (.A1(_02374_),
    .A2(_02383_),
    .B1(_02408_),
    .Y(_02410_));
 sky130_fd_sc_hd__nor3_2 _11616_ (.A(_02404_),
    .B(_02409_),
    .C(_02410_),
    .Y(_02411_));
 sky130_fd_sc_hd__or3_2 _11617_ (.A(_02404_),
    .B(_02409_),
    .C(_02410_),
    .X(_02412_));
 sky130_fd_sc_hd__o211ai_4 _11618_ (.A1(_02409_),
    .A2(_02411_),
    .B1(_02377_),
    .C1(_02382_),
    .Y(_02413_));
 sky130_fd_sc_hd__o21ba_1 _11619_ (.A1(_02336_),
    .A2(_02345_),
    .B1_N(_02378_),
    .X(_02414_));
 sky130_fd_sc_hd__nor3_1 _11620_ (.A(_02379_),
    .B(_02413_),
    .C(_02414_),
    .Y(_02415_));
 sky130_fd_sc_hd__o21a_1 _11621_ (.A1(_02379_),
    .A2(_02414_),
    .B1(_02413_),
    .X(_02416_));
 sky130_fd_sc_hd__or2_1 _11622_ (.A(_02415_),
    .B(_02416_),
    .X(_02417_));
 sky130_fd_sc_hd__a211o_1 _11623_ (.A1(_02377_),
    .A2(_02382_),
    .B1(_02409_),
    .C1(_02411_),
    .X(_02418_));
 sky130_fd_sc_hd__nand2_1 _11624_ (.A(_02413_),
    .B(_02418_),
    .Y(_02419_));
 sky130_fd_sc_hd__o21ai_2 _11625_ (.A1(_02409_),
    .A2(_02410_),
    .B1(_02404_),
    .Y(_02420_));
 sky130_fd_sc_hd__and2_1 _11626_ (.A(_02412_),
    .B(_02420_),
    .X(_02421_));
 sky130_fd_sc_hd__a21o_1 _11627_ (.A1(_02402_),
    .A2(_02403_),
    .B1(_02406_),
    .X(_02422_));
 sky130_fd_sc_hd__xnor2_4 _11628_ (.A(_02389_),
    .B(_02390_),
    .Y(_02423_));
 sky130_fd_sc_hd__and4_1 _11629_ (.A(net591),
    .B(net614),
    .C(net889),
    .D(net905),
    .X(_02424_));
 sky130_fd_sc_hd__nand2_4 _11630_ (.A(net603),
    .B(net899),
    .Y(_02425_));
 sky130_fd_sc_hd__a22oi_2 _11631_ (.A1(net614),
    .A2(net889),
    .B1(net905),
    .B2(net591),
    .Y(_02426_));
 sky130_fd_sc_hd__or2_4 _11632_ (.A(_02424_),
    .B(_02426_),
    .X(_02427_));
 sky130_fd_sc_hd__o21ba_2 _11633_ (.A1(_02425_),
    .A2(_02426_),
    .B1_N(_02424_),
    .X(_02428_));
 sky130_fd_sc_hd__nand2b_1 _11634_ (.A_N(_02428_),
    .B(_02423_),
    .Y(_02429_));
 sky130_fd_sc_hd__xnor2_4 _11635_ (.A(_02423_),
    .B(_02428_),
    .Y(_02430_));
 sky130_fd_sc_hd__o22a_1 _11636_ (.A1(net304),
    .A2(net282),
    .B1(_03302_),
    .B2(net309),
    .X(_02431_));
 sky130_fd_sc_hd__nor2_2 _11637_ (.A(_02348_),
    .B(_02431_),
    .Y(_02432_));
 sky130_fd_sc_hd__nand2_2 _11638_ (.A(_02430_),
    .B(_02432_),
    .Y(_02433_));
 sky130_fd_sc_hd__xnor2_2 _11639_ (.A(_02393_),
    .B(_02395_),
    .Y(_02434_));
 sky130_fd_sc_hd__nor2_4 _11640_ (.A(_02433_),
    .B(_02434_),
    .Y(_02435_));
 sky130_fd_sc_hd__xor2_4 _11641_ (.A(_02392_),
    .B(_02435_),
    .X(_02436_));
 sky130_fd_sc_hd__a22o_1 _11642_ (.A1(net533),
    .A2(net917),
    .B1(_02398_),
    .B2(_02399_),
    .X(_02437_));
 sky130_fd_sc_hd__nand2b_1 _11643_ (.A_N(_02400_),
    .B(_02437_),
    .Y(_02438_));
 sky130_fd_sc_hd__and3b_1 _11644_ (.A_N(_02400_),
    .B(_02436_),
    .C(_02437_),
    .X(_02439_));
 sky130_fd_sc_hd__a21o_1 _11645_ (.A1(_02392_),
    .A2(_02435_),
    .B1(_02439_),
    .X(_02440_));
 sky130_fd_sc_hd__and3_2 _11646_ (.A(_02407_),
    .B(_02422_),
    .C(_02440_),
    .X(_02441_));
 sky130_fd_sc_hd__a22o_1 _11647_ (.A1(_02413_),
    .A2(_02418_),
    .B1(_02421_),
    .B2(_02441_),
    .X(_02442_));
 sky130_fd_sc_hd__xnor2_2 _11648_ (.A(_02436_),
    .B(_02438_),
    .Y(_02443_));
 sky130_fd_sc_hd__xor2_4 _11649_ (.A(_02425_),
    .B(_02427_),
    .X(_02444_));
 sky130_fd_sc_hd__a22o_1 _11650_ (.A1(net615),
    .A2(net899),
    .B1(net914),
    .B2(net591),
    .X(_02445_));
 sky130_fd_sc_hd__nand2_4 _11651_ (.A(net615),
    .B(net914),
    .Y(_02446_));
 sky130_fd_sc_hd__nor2_2 _11652_ (.A(_02387_),
    .B(_02446_),
    .Y(_02447_));
 sky130_fd_sc_hd__nor2_2 _11653_ (.A(net292),
    .B(net282),
    .Y(_02448_));
 sky130_fd_sc_hd__o21a_1 _11654_ (.A1(_02387_),
    .A2(_02446_),
    .B1(_02445_),
    .X(_02449_));
 sky130_fd_sc_hd__and2_1 _11655_ (.A(_02448_),
    .B(_02449_),
    .X(_02450_));
 sky130_fd_sc_hd__o21ai_4 _11656_ (.A1(_02447_),
    .A2(_02450_),
    .B1(_02444_),
    .Y(_02451_));
 sky130_fd_sc_hd__or3_2 _11657_ (.A(_02444_),
    .B(_02447_),
    .C(_02450_),
    .X(_02452_));
 sky130_fd_sc_hd__nand4_2 _11658_ (.A(net579),
    .B(net915),
    .C(_02451_),
    .D(_02452_),
    .Y(_02453_));
 sky130_fd_sc_hd__xnor2_2 _11659_ (.A(_02430_),
    .B(_02432_),
    .Y(_02454_));
 sky130_fd_sc_hd__nor2_1 _11660_ (.A(_02453_),
    .B(_02454_),
    .Y(_02455_));
 sky130_fd_sc_hd__and2b_1 _11661_ (.A_N(_02429_),
    .B(_02455_),
    .X(_02456_));
 sky130_fd_sc_hd__xnor2_1 _11662_ (.A(_02429_),
    .B(_02455_),
    .Y(_02457_));
 sky130_fd_sc_hd__and2_1 _11663_ (.A(_02433_),
    .B(_02434_),
    .X(_02458_));
 sky130_fd_sc_hd__nor2_1 _11664_ (.A(_02435_),
    .B(_02458_),
    .Y(_02459_));
 sky130_fd_sc_hd__and2_1 _11665_ (.A(_02457_),
    .B(_02459_),
    .X(_02460_));
 sky130_fd_sc_hd__nor2_2 _11666_ (.A(_02456_),
    .B(_02460_),
    .Y(_02461_));
 sky130_fd_sc_hd__and2b_1 _11667_ (.A_N(_02461_),
    .B(_02443_),
    .X(_02462_));
 sky130_fd_sc_hd__a21o_1 _11668_ (.A1(_02407_),
    .A2(_02422_),
    .B1(_02440_),
    .X(_02463_));
 sky130_fd_sc_hd__and2b_1 _11669_ (.A_N(_02441_),
    .B(_02463_),
    .X(_02464_));
 sky130_fd_sc_hd__and3b_1 _11670_ (.A_N(_02441_),
    .B(_02462_),
    .C(_02463_),
    .X(_02465_));
 sky130_fd_sc_hd__or2_1 _11671_ (.A(_02441_),
    .B(_02465_),
    .X(_02466_));
 sky130_fd_sc_hd__nand3_2 _11672_ (.A(_02412_),
    .B(_02420_),
    .C(_02466_),
    .Y(_02467_));
 sky130_fd_sc_hd__nor2_1 _11673_ (.A(_02457_),
    .B(_02459_),
    .Y(_02468_));
 sky130_fd_sc_hd__or2_2 _11674_ (.A(_02460_),
    .B(_02468_),
    .X(_02469_));
 sky130_fd_sc_hd__or3_1 _11675_ (.A(net292),
    .B(net282),
    .C(_02446_),
    .X(_02470_));
 sky130_fd_sc_hd__nor2_1 _11676_ (.A(_02449_),
    .B(_02470_),
    .Y(_02471_));
 sky130_fd_sc_hd__a22o_1 _11677_ (.A1(net579),
    .A2(net915),
    .B1(_02451_),
    .B2(_02452_),
    .X(_02472_));
 sky130_fd_sc_hd__and2_1 _11678_ (.A(_02453_),
    .B(_02472_),
    .X(_02473_));
 sky130_fd_sc_hd__nand2_1 _11679_ (.A(_02471_),
    .B(_02473_),
    .Y(_02474_));
 sky130_fd_sc_hd__nor2_1 _11680_ (.A(_02451_),
    .B(_02454_),
    .Y(_02475_));
 sky130_fd_sc_hd__or2_2 _11681_ (.A(_02451_),
    .B(_02454_),
    .X(_02476_));
 sky130_fd_sc_hd__a311o_1 _11682_ (.A1(_02451_),
    .A2(_02453_),
    .A3(_02454_),
    .B1(_02455_),
    .C1(_02475_),
    .X(_02477_));
 sky130_fd_sc_hd__or2_2 _11683_ (.A(_02474_),
    .B(_02477_),
    .X(_02478_));
 sky130_fd_sc_hd__nor2_1 _11684_ (.A(_02469_),
    .B(_02478_),
    .Y(_02479_));
 sky130_fd_sc_hd__nor2_1 _11685_ (.A(_02469_),
    .B(_02476_),
    .Y(_02480_));
 sky130_fd_sc_hd__xnor2_2 _11686_ (.A(_02443_),
    .B(_02461_),
    .Y(_02481_));
 sky130_fd_sc_hd__nand2_1 _11687_ (.A(_02480_),
    .B(_02481_),
    .Y(_02482_));
 sky130_fd_sc_hd__xor2_1 _11688_ (.A(_02480_),
    .B(_02481_),
    .X(_02483_));
 sky130_fd_sc_hd__nand2_1 _11689_ (.A(_02479_),
    .B(_02483_),
    .Y(_02484_));
 sky130_fd_sc_hd__xnor2_1 _11690_ (.A(_02462_),
    .B(_02464_),
    .Y(_02485_));
 sky130_fd_sc_hd__nor2_1 _11691_ (.A(_02484_),
    .B(_02485_),
    .Y(_02486_));
 sky130_fd_sc_hd__or3b_1 _11692_ (.A(_02441_),
    .B(_02482_),
    .C_N(_02463_),
    .X(_02487_));
 sky130_fd_sc_hd__inv_2 _11693_ (.A(_02487_),
    .Y(_02488_));
 sky130_fd_sc_hd__a21o_1 _11694_ (.A1(_02412_),
    .A2(_02420_),
    .B1(_02466_),
    .X(_02489_));
 sky130_fd_sc_hd__o211a_1 _11695_ (.A1(_02486_),
    .A2(_02488_),
    .B1(_02489_),
    .C1(_02467_),
    .X(_02490_));
 sky130_fd_sc_hd__o2bb2a_2 _11696_ (.A1_N(_02442_),
    .A2_N(_02490_),
    .B1(_02467_),
    .B2(_02419_),
    .X(_02491_));
 sky130_fd_sc_hd__nor2_1 _11697_ (.A(_02417_),
    .B(_02491_),
    .Y(_02492_));
 sky130_fd_sc_hd__o21bai_2 _11698_ (.A1(_02416_),
    .A2(_02491_),
    .B1_N(_02415_),
    .Y(_02493_));
 sky130_fd_sc_hd__a21o_1 _11699_ (.A1(_02338_),
    .A2(_02380_),
    .B1(_02379_),
    .X(_02494_));
 sky130_fd_sc_hd__nand3_1 _11700_ (.A(_02381_),
    .B(_02493_),
    .C(_02494_),
    .Y(_02495_));
 sky130_fd_sc_hd__a21bo_1 _11701_ (.A1(_02493_),
    .A2(_02494_),
    .B1_N(_02381_),
    .X(_02496_));
 sky130_fd_sc_hd__nand2_1 _11702_ (.A(_02344_),
    .B(_02496_),
    .Y(_02497_));
 sky130_fd_sc_hd__xor2_4 _11703_ (.A(_02214_),
    .B(_02256_),
    .X(_02498_));
 sky130_fd_sc_hd__xnor2_4 _11704_ (.A(_02340_),
    .B(_02498_),
    .Y(_02499_));
 sky130_fd_sc_hd__nand2_1 _11705_ (.A(_02340_),
    .B(_02342_),
    .Y(_02500_));
 sky130_fd_sc_hd__a32o_2 _11706_ (.A1(_02344_),
    .A2(_02496_),
    .A3(_02499_),
    .B1(_02500_),
    .B2(_02498_),
    .X(_02501_));
 sky130_fd_sc_hd__nand2_2 _11707_ (.A(_02260_),
    .B(_02501_),
    .Y(_02502_));
 sky130_fd_sc_hd__xor2_4 _11708_ (.A(_02208_),
    .B(_02213_),
    .X(_02503_));
 sky130_fd_sc_hd__o21bai_1 _11709_ (.A1(_02257_),
    .A2(_02258_),
    .B1_N(_02208_),
    .Y(_02504_));
 sky130_fd_sc_hd__a32o_2 _11710_ (.A1(_02260_),
    .A2(_02501_),
    .A3(_02503_),
    .B1(_02504_),
    .B2(_02213_),
    .X(_02505_));
 sky130_fd_sc_hd__xnor2_4 _11711_ (.A(_02029_),
    .B(_02095_),
    .Y(_02506_));
 sky130_fd_sc_hd__and2_1 _11712_ (.A(_02212_),
    .B(_02506_),
    .X(_02507_));
 sky130_fd_sc_hd__xor2_4 _11713_ (.A(_02212_),
    .B(_02506_),
    .X(_02508_));
 sky130_fd_sc_hd__and2_1 _11714_ (.A(_02505_),
    .B(_02508_),
    .X(_02509_));
 sky130_fd_sc_hd__and3_2 _11715_ (.A(_02097_),
    .B(_02505_),
    .C(_02508_),
    .X(_02510_));
 sky130_fd_sc_hd__o21a_2 _11716_ (.A1(_02096_),
    .A2(_02507_),
    .B1(_02027_),
    .X(_02511_));
 sky130_fd_sc_hd__and3_1 _11717_ (.A(_02025_),
    .B(_02097_),
    .C(_02508_),
    .X(_02512_));
 sky130_fd_sc_hd__a221o_4 _11718_ (.A1(_02025_),
    .A2(_02511_),
    .B1(_02512_),
    .B2(_02505_),
    .C1(_02026_),
    .X(_02513_));
 sky130_fd_sc_hd__and2_2 _11719_ (.A(_02002_),
    .B(_02004_),
    .X(_02514_));
 sky130_fd_sc_hd__or2_4 _11720_ (.A(_01552_),
    .B(_02514_),
    .X(_02515_));
 sky130_fd_sc_hd__o21a_1 _11721_ (.A1(_01562_),
    .A2(_01568_),
    .B1(_01567_),
    .X(_02516_));
 sky130_fd_sc_hd__nor2_2 _11722_ (.A(_01569_),
    .B(_02516_),
    .Y(_02517_));
 sky130_fd_sc_hd__a21bo_2 _11723_ (.A1(_01526_),
    .A2(_01560_),
    .B1_N(_01559_),
    .X(_02518_));
 sky130_fd_sc_hd__o21ai_4 _11724_ (.A1(_02006_),
    .A2(_02010_),
    .B1(_02009_),
    .Y(_02519_));
 sky130_fd_sc_hd__and3_4 _11725_ (.A(_01561_),
    .B(_02518_),
    .C(_02519_),
    .X(_02520_));
 sky130_fd_sc_hd__nand2_1 _11726_ (.A(_01552_),
    .B(_02514_),
    .Y(_02521_));
 sky130_fd_sc_hd__nand2_2 _11727_ (.A(_02515_),
    .B(_02521_),
    .Y(_02522_));
 sky130_fd_sc_hd__a21oi_4 _11728_ (.A1(_01561_),
    .A2(_02518_),
    .B1(_02519_),
    .Y(_02523_));
 sky130_fd_sc_hd__nor3_4 _11729_ (.A(_02520_),
    .B(_02522_),
    .C(_02523_),
    .Y(_02524_));
 sky130_fd_sc_hd__o21a_2 _11730_ (.A1(_02520_),
    .A2(_02524_),
    .B1(_02517_),
    .X(_02525_));
 sky130_fd_sc_hd__nor3_4 _11731_ (.A(_02517_),
    .B(_02520_),
    .C(_02524_),
    .Y(_02526_));
 sky130_fd_sc_hd__nor3_4 _11732_ (.A(_02515_),
    .B(_02525_),
    .C(_02526_),
    .Y(_02527_));
 sky130_fd_sc_hd__o21a_2 _11733_ (.A1(_02525_),
    .A2(_02526_),
    .B1(_02515_),
    .X(_02528_));
 sky130_fd_sc_hd__o21a_1 _11734_ (.A1(_02520_),
    .A2(_02523_),
    .B1(_02522_),
    .X(_02529_));
 sky130_fd_sc_hd__o21ai_1 _11735_ (.A1(_02000_),
    .A2(_02015_),
    .B1(_02014_),
    .Y(_02530_));
 sky130_fd_sc_hd__nor3b_2 _11736_ (.A(_02524_),
    .B(_02529_),
    .C_N(_02530_),
    .Y(_02531_));
 sky130_fd_sc_hd__inv_2 _11737_ (.A(_02531_),
    .Y(_02532_));
 sky130_fd_sc_hd__o21ba_1 _11738_ (.A1(_02524_),
    .A2(_02529_),
    .B1_N(_02530_),
    .X(_02533_));
 sky130_fd_sc_hd__or3_4 _11739_ (.A(_01998_),
    .B(_02531_),
    .C(_02533_),
    .X(_02534_));
 sky130_fd_sc_hd__a211oi_4 _11740_ (.A1(_02532_),
    .A2(_02534_),
    .B1(_02527_),
    .C1(_02528_),
    .Y(_02535_));
 sky130_fd_sc_hd__o21a_1 _11741_ (.A1(_01570_),
    .A2(_01571_),
    .B1(_01565_),
    .X(_02536_));
 sky130_fd_sc_hd__or2_2 _11742_ (.A(_01572_),
    .B(_02536_),
    .X(_02537_));
 sky130_fd_sc_hd__o21bai_4 _11743_ (.A1(_02515_),
    .A2(_02526_),
    .B1_N(_02525_),
    .Y(_02538_));
 sky130_fd_sc_hd__nand2b_4 _11744_ (.A_N(_02537_),
    .B(_02538_),
    .Y(_02539_));
 sky130_fd_sc_hd__xnor2_1 _11745_ (.A(_02537_),
    .B(_02538_),
    .Y(_02540_));
 sky130_fd_sc_hd__nand2_1 _11746_ (.A(_02535_),
    .B(_02540_),
    .Y(_02541_));
 sky130_fd_sc_hd__or2_1 _11747_ (.A(_02535_),
    .B(_02540_),
    .X(_02542_));
 sky130_fd_sc_hd__and2_2 _11748_ (.A(_02541_),
    .B(_02542_),
    .X(_02543_));
 sky130_fd_sc_hd__xnor2_4 _11749_ (.A(_01355_),
    .B(_01574_),
    .Y(_02544_));
 sky130_fd_sc_hd__xor2_4 _11750_ (.A(_02539_),
    .B(_02544_),
    .X(_02545_));
 sky130_fd_sc_hd__o21ai_1 _11751_ (.A1(_02531_),
    .A2(_02533_),
    .B1(_01998_),
    .Y(_02546_));
 sky130_fd_sc_hd__a21o_1 _11752_ (.A1(_02016_),
    .A2(_02017_),
    .B1(_02019_),
    .X(_02547_));
 sky130_fd_sc_hd__and3_4 _11753_ (.A(_02534_),
    .B(_02546_),
    .C(_02547_),
    .X(_02548_));
 sky130_fd_sc_hd__a21o_1 _11754_ (.A1(_02534_),
    .A2(_02546_),
    .B1(_02547_),
    .X(_02549_));
 sky130_fd_sc_hd__and2b_2 _11755_ (.A_N(_02548_),
    .B(_02549_),
    .X(_02550_));
 sky130_fd_sc_hd__xor2_4 _11756_ (.A(_02022_),
    .B(_02550_),
    .X(_02551_));
 sky130_fd_sc_hd__o211a_1 _11757_ (.A1(_02527_),
    .A2(_02528_),
    .B1(_02532_),
    .C1(_02534_),
    .X(_02552_));
 sky130_fd_sc_hd__nor2_4 _11758_ (.A(_02535_),
    .B(_02552_),
    .Y(_02553_));
 sky130_fd_sc_hd__xor2_4 _11759_ (.A(_02548_),
    .B(_02553_),
    .X(_02554_));
 sky130_fd_sc_hd__and4_1 _11760_ (.A(_02543_),
    .B(_02545_),
    .C(_02551_),
    .D(_02554_),
    .X(_02555_));
 sky130_fd_sc_hd__a21o_1 _11761_ (.A1(_02022_),
    .A2(_02549_),
    .B1(_02548_),
    .X(_02556_));
 sky130_fd_sc_hd__and2_1 _11762_ (.A(_02553_),
    .B(_02556_),
    .X(_02557_));
 sky130_fd_sc_hd__a21oi_1 _11763_ (.A1(_02539_),
    .A2(_02541_),
    .B1(_02544_),
    .Y(_02558_));
 sky130_fd_sc_hd__a31o_1 _11764_ (.A1(_02543_),
    .A2(_02545_),
    .A3(_02557_),
    .B1(_02558_),
    .X(_02559_));
 sky130_fd_sc_hd__a21oi_4 _11765_ (.A1(_02513_),
    .A2(_02555_),
    .B1(_02559_),
    .Y(_02560_));
 sky130_fd_sc_hd__or2_1 _11766_ (.A(_01579_),
    .B(_02560_),
    .X(_02561_));
 sky130_fd_sc_hd__or2_2 _11767_ (.A(_01481_),
    .B(_01578_),
    .X(_02562_));
 sky130_fd_sc_hd__or2_1 _11768_ (.A(_01481_),
    .B(_01577_),
    .X(_02563_));
 sky130_fd_sc_hd__o31ai_4 _11769_ (.A1(_01481_),
    .A2(_01579_),
    .A3(_02560_),
    .B1(_02562_),
    .Y(_02564_));
 sky130_fd_sc_hd__a21boi_1 _11770_ (.A1(_01375_),
    .A2(_01376_),
    .B1_N(_01263_),
    .Y(_02565_));
 sky130_fd_sc_hd__nand2_1 _11771_ (.A(_01263_),
    .B(_01376_),
    .Y(_02566_));
 sky130_fd_sc_hd__a31o_1 _11772_ (.A1(_01263_),
    .A2(_01378_),
    .A3(_02564_),
    .B1(_02565_),
    .X(_02567_));
 sky130_fd_sc_hd__and2_1 _11773_ (.A(_01145_),
    .B(_02567_),
    .X(_02568_));
 sky130_fd_sc_hd__a21boi_1 _11774_ (.A1(_01142_),
    .A2(_01143_),
    .B1_N(_01020_),
    .Y(_02569_));
 sky130_fd_sc_hd__nand2_1 _11775_ (.A(_01020_),
    .B(_01143_),
    .Y(_02570_));
 sky130_fd_sc_hd__a31o_4 _11776_ (.A1(_01020_),
    .A2(_01145_),
    .A3(_02567_),
    .B1(_02569_),
    .X(_02571_));
 sky130_fd_sc_hd__a21boi_1 _11777_ (.A1(_00890_),
    .A2(_00891_),
    .B1_N(_00763_),
    .Y(_02572_));
 sky130_fd_sc_hd__nand2_2 _11778_ (.A(_00763_),
    .B(_00891_),
    .Y(_02573_));
 sky130_fd_sc_hd__a31o_4 _11779_ (.A1(_00763_),
    .A2(_00893_),
    .A3(_02571_),
    .B1(_02572_),
    .X(_02574_));
 sky130_fd_sc_hd__inv_2 _11780_ (.A(_02574_),
    .Y(_02575_));
 sky130_fd_sc_hd__and2_1 _11781_ (.A(_00621_),
    .B(_02574_),
    .X(_02576_));
 sky130_fd_sc_hd__nand2b_4 _11782_ (.A_N(net316),
    .B(net315),
    .Y(_02577_));
 sky130_fd_sc_hd__nor2_2 _11783_ (.A(_03452_),
    .B(_02577_),
    .Y(_02578_));
 sky130_fd_sc_hd__or2_2 _11784_ (.A(_03452_),
    .B(_02577_),
    .X(_02579_));
 sky130_fd_sc_hd__o21a_1 _11785_ (.A1(_00619_),
    .A2(_02576_),
    .B1(_00474_),
    .X(_02580_));
 sky130_fd_sc_hd__o31ai_2 _11786_ (.A1(_00474_),
    .A2(_00619_),
    .A3(_02576_),
    .B1(net260),
    .Y(_02581_));
 sky130_fd_sc_hd__or2_4 _11787_ (.A(net515),
    .B(net523),
    .X(_02582_));
 sky130_fd_sc_hd__or2_4 _11788_ (.A(net451),
    .B(net461),
    .X(_02583_));
 sky130_fd_sc_hd__or3_4 _11789_ (.A(net451),
    .B(net461),
    .C(net471),
    .X(_02584_));
 sky130_fd_sc_hd__or2_1 _11790_ (.A(net471),
    .B(net478),
    .X(_02585_));
 sky130_fd_sc_hd__or4_2 _11791_ (.A(net451),
    .B(net461),
    .C(net471),
    .D(net478),
    .X(_02586_));
 sky130_fd_sc_hd__or3_4 _11792_ (.A(net471),
    .B(net478),
    .C(net490),
    .X(_02587_));
 sky130_fd_sc_hd__or2_2 _11793_ (.A(net500),
    .B(net507),
    .X(_02588_));
 sky130_fd_sc_hd__or4_1 _11794_ (.A(net386),
    .B(net395),
    .C(net402),
    .D(net410),
    .X(_02589_));
 sky130_fd_sc_hd__or4_1 _11795_ (.A(net417),
    .B(net426),
    .C(net434),
    .D(net444),
    .X(_02590_));
 sky130_fd_sc_hd__or4_1 _11796_ (.A(net354),
    .B(net361),
    .C(net370),
    .D(net379),
    .X(_02591_));
 sky130_fd_sc_hd__or4_1 _11797_ (.A(net319),
    .B(net330),
    .C(net336),
    .D(net348),
    .X(_02592_));
 sky130_fd_sc_hd__or4_4 _11798_ (.A(_02583_),
    .B(_02589_),
    .C(_02591_),
    .D(_02592_),
    .X(_02593_));
 sky130_fd_sc_hd__or2_2 _11799_ (.A(_02587_),
    .B(_02590_),
    .X(_02594_));
 sky130_fd_sc_hd__nor4_4 _11800_ (.A(_02582_),
    .B(_02588_),
    .C(_02593_),
    .D(_02594_),
    .Y(_02595_));
 sky130_fd_sc_hd__a21o_1 _11801_ (.A1(net284),
    .A2(net724),
    .B1(_01337_),
    .X(_02596_));
 sky130_fd_sc_hd__nand2_1 _11802_ (.A(net213),
    .B(_02596_),
    .Y(_02597_));
 sky130_fd_sc_hd__a21o_1 _11803_ (.A1(net283),
    .A2(net704),
    .B1(_01103_),
    .X(_02598_));
 sky130_fd_sc_hd__nand2_1 _11804_ (.A(net213),
    .B(_02598_),
    .Y(_02599_));
 sky130_fd_sc_hd__mux2_1 _11805_ (.A0(_02597_),
    .A1(_02599_),
    .S(net287),
    .X(_02600_));
 sky130_fd_sc_hd__a21o_1 _11806_ (.A1(net283),
    .A2(net687),
    .B1(_00720_),
    .X(_02601_));
 sky130_fd_sc_hd__nand2_1 _11807_ (.A(net213),
    .B(_02601_),
    .Y(_02602_));
 sky130_fd_sc_hd__and2_1 _11808_ (.A(net283),
    .B(net669),
    .X(_02603_));
 sky130_fd_sc_hd__o21ai_2 _11809_ (.A1(_00446_),
    .A2(_02603_),
    .B1(net212),
    .Y(_02604_));
 sky130_fd_sc_hd__mux2_1 _11810_ (.A0(_02602_),
    .A1(_02604_),
    .S(net288),
    .X(_02605_));
 sky130_fd_sc_hd__and2_1 _11811_ (.A(net283),
    .B(net618),
    .X(_02606_));
 sky130_fd_sc_hd__o21a_1 _11812_ (.A1(_07313_),
    .A2(_02606_),
    .B1(net212),
    .X(_02607_));
 sky130_fd_sc_hd__and2_1 _11813_ (.A(net283),
    .B(net653),
    .X(_02608_));
 sky130_fd_sc_hd__o21ai_1 _11814_ (.A1(_00144_),
    .A2(_02608_),
    .B1(net212),
    .Y(_02609_));
 sky130_fd_sc_hd__and2_1 _11815_ (.A(net283),
    .B(\cla_inst.in1[29] ),
    .X(_02610_));
 sky130_fd_sc_hd__o21ai_1 _11816_ (.A1(_07302_),
    .A2(_02610_),
    .B1(net212),
    .Y(_02611_));
 sky130_fd_sc_hd__mux2_1 _11817_ (.A0(_02609_),
    .A1(_02611_),
    .S(net287),
    .X(_02612_));
 sky130_fd_sc_hd__nor2_1 _11818_ (.A(net293),
    .B(_02612_),
    .Y(_02613_));
 sky130_fd_sc_hd__a31o_2 _11819_ (.A1(net293),
    .A2(net598),
    .A3(_02607_),
    .B1(_02613_),
    .X(_02614_));
 sky130_fd_sc_hd__inv_2 _11820_ (.A(_02614_),
    .Y(_02615_));
 sky130_fd_sc_hd__mux4_1 _11821_ (.A0(_02597_),
    .A1(_02599_),
    .A2(_02602_),
    .A3(_02604_),
    .S0(net287),
    .S1(net294),
    .X(_02616_));
 sky130_fd_sc_hd__mux2_1 _11822_ (.A0(_02615_),
    .A1(_02616_),
    .S(net566),
    .X(_02617_));
 sky130_fd_sc_hd__mux2_1 _11823_ (.A0(net891),
    .A1(net900),
    .S(net608),
    .X(_02618_));
 sky130_fd_sc_hd__nand2_1 _11824_ (.A(net215),
    .B(_02618_),
    .Y(_02619_));
 sky130_fd_sc_hd__a21bo_1 _11825_ (.A1(net286),
    .A2(net865),
    .B1_N(_02312_),
    .X(_02620_));
 sky130_fd_sc_hd__nand2_2 _11826_ (.A(_02595_),
    .B(_02620_),
    .Y(_02621_));
 sky130_fd_sc_hd__mux2_1 _11827_ (.A0(_02619_),
    .A1(_02621_),
    .S(net288),
    .X(_02622_));
 sky130_fd_sc_hd__mux2_1 _11828_ (.A0(net842),
    .A1(\ApproximateM_inst.lob_16.lob1.genblk1[6].genblk1.mux.sel ),
    .S(net606),
    .X(_02623_));
 sky130_fd_sc_hd__nand2_1 _11829_ (.A(net212),
    .B(_02623_),
    .Y(_02624_));
 sky130_fd_sc_hd__mux2_1 _11830_ (.A0(net823),
    .A1(net832),
    .S(net606),
    .X(_02625_));
 sky130_fd_sc_hd__nand2_1 _11831_ (.A(net212),
    .B(_02625_),
    .Y(_02626_));
 sky130_fd_sc_hd__mux2_1 _11832_ (.A0(_02624_),
    .A1(_02626_),
    .S(net288),
    .X(_02627_));
 sky130_fd_sc_hd__mux2_1 _11833_ (.A0(_02622_),
    .A1(_02627_),
    .S(net293),
    .X(_02628_));
 sky130_fd_sc_hd__mux2_1 _11834_ (.A0(net803),
    .A1(net813),
    .S(net606),
    .X(_02629_));
 sky130_fd_sc_hd__nand2_1 _11835_ (.A(net212),
    .B(_02629_),
    .Y(_02630_));
 sky130_fd_sc_hd__mux2_1 _11836_ (.A0(net777),
    .A1(net788),
    .S(net606),
    .X(_02631_));
 sky130_fd_sc_hd__nand2_1 _11837_ (.A(net212),
    .B(_02631_),
    .Y(_02632_));
 sky130_fd_sc_hd__mux2_1 _11838_ (.A0(_02630_),
    .A1(_02632_),
    .S(net287),
    .X(_02633_));
 sky130_fd_sc_hd__mux2_1 _11839_ (.A0(net760),
    .A1(net771),
    .S(net606),
    .X(_02634_));
 sky130_fd_sc_hd__nand2_1 _11840_ (.A(net212),
    .B(_02634_),
    .Y(_02635_));
 sky130_fd_sc_hd__and2_2 _11841_ (.A(net286),
    .B(net745),
    .X(_02636_));
 sky130_fd_sc_hd__o21ai_4 _11842_ (.A1(_01547_),
    .A2(_02636_),
    .B1(net217),
    .Y(_02637_));
 sky130_fd_sc_hd__mux2_1 _11843_ (.A0(_02635_),
    .A1(_02637_),
    .S(net287),
    .X(_02638_));
 sky130_fd_sc_hd__mux4_2 _11844_ (.A0(_02622_),
    .A1(_02627_),
    .A2(_02633_),
    .A3(_02638_),
    .S0(net294),
    .S1(net302),
    .X(_02639_));
 sky130_fd_sc_hd__mux2_1 _11845_ (.A0(_02617_),
    .A1(_02639_),
    .S(net552),
    .X(_02640_));
 sky130_fd_sc_hd__nor3_4 _11846_ (.A(net534),
    .B(_03420_),
    .C(_02577_),
    .Y(_02641_));
 sky130_fd_sc_hd__or3_4 _11847_ (.A(net534),
    .B(_03420_),
    .C(_02577_),
    .X(_02642_));
 sky130_fd_sc_hd__nor2_2 _11848_ (.A(net537),
    .B(_02642_),
    .Y(_02643_));
 sky130_fd_sc_hd__nand2_2 _11849_ (.A(_03193_),
    .B(_02641_),
    .Y(_02644_));
 sky130_fd_sc_hd__o21ai_1 _11850_ (.A1(net611),
    .A2(net282),
    .B1(_02446_),
    .Y(_02645_));
 sky130_fd_sc_hd__nand2_2 _11851_ (.A(net216),
    .B(_02645_),
    .Y(_02646_));
 sky130_fd_sc_hd__or2_2 _11852_ (.A(net597),
    .B(_02646_),
    .X(_02647_));
 sky130_fd_sc_hd__nand2_2 _11853_ (.A(net308),
    .B(_02641_),
    .Y(_02648_));
 sky130_fd_sc_hd__or3_4 _11854_ (.A(net566),
    .B(net584),
    .C(_02647_),
    .X(_02649_));
 sky130_fd_sc_hd__o21a_1 _11855_ (.A1(net552),
    .A2(_02649_),
    .B1(net540),
    .X(_02650_));
 sky130_fd_sc_hd__a211o_2 _11856_ (.A1(_03193_),
    .A2(_02640_),
    .B1(_02642_),
    .C1(_02650_),
    .X(_02651_));
 sky130_fd_sc_hd__o21ai_2 _11857_ (.A1(_02580_),
    .A2(_02581_),
    .B1(_02651_),
    .Y(_08653_));
 sky130_fd_sc_hd__a22oi_4 _11858_ (.A1(net421),
    .A2(net746),
    .B1(net767),
    .B2(net404),
    .Y(_02652_));
 sky130_fd_sc_hd__and4_1 _11859_ (.A(net404),
    .B(net421),
    .C(net747),
    .D(net767),
    .X(_02653_));
 sky130_fd_sc_hd__nor2_2 _11860_ (.A(_02652_),
    .B(_02653_),
    .Y(_02654_));
 sky130_fd_sc_hd__nand2_4 _11861_ (.A(net413),
    .B(net756),
    .Y(_02655_));
 sky130_fd_sc_hd__xnor2_4 _11862_ (.A(_02654_),
    .B(_02655_),
    .Y(_02656_));
 sky130_fd_sc_hd__a31o_2 _11863_ (.A1(net413),
    .A2(net767),
    .A3(_03484_),
    .B1(_03495_),
    .X(_02657_));
 sky130_fd_sc_hd__nand2_2 _11864_ (.A(_02656_),
    .B(_02657_),
    .Y(_02658_));
 sky130_fd_sc_hd__xor2_2 _11865_ (.A(_02656_),
    .B(_02657_),
    .X(_02659_));
 sky130_fd_sc_hd__a22oi_1 _11866_ (.A1(net436),
    .A2(net730),
    .B1(net738),
    .B2(net428),
    .Y(_02660_));
 sky130_fd_sc_hd__and4_2 _11867_ (.A(net428),
    .B(net436),
    .C(net730),
    .D(net738),
    .X(_02661_));
 sky130_fd_sc_hd__nor2_1 _11868_ (.A(_02660_),
    .B(_02661_),
    .Y(_02662_));
 sky130_fd_sc_hd__nand2_1 _11869_ (.A(net446),
    .B(net721),
    .Y(_02663_));
 sky130_fd_sc_hd__and3_2 _11870_ (.A(net446),
    .B(net721),
    .C(_02662_),
    .X(_02664_));
 sky130_fd_sc_hd__xor2_1 _11871_ (.A(_02662_),
    .B(_02663_),
    .X(_02665_));
 sky130_fd_sc_hd__inv_2 _11872_ (.A(_02665_),
    .Y(_02666_));
 sky130_fd_sc_hd__nand2_2 _11873_ (.A(_02659_),
    .B(_02666_),
    .Y(_02667_));
 sky130_fd_sc_hd__or2_1 _11874_ (.A(_02659_),
    .B(_02666_),
    .X(_02668_));
 sky130_fd_sc_hd__nand2_2 _11875_ (.A(_02667_),
    .B(_02668_),
    .Y(_02669_));
 sky130_fd_sc_hd__a21oi_4 _11876_ (.A1(_03604_),
    .A2(_03702_),
    .B1(_02669_),
    .Y(_02670_));
 sky130_fd_sc_hd__and3_2 _11877_ (.A(_03604_),
    .B(_03702_),
    .C(_02669_),
    .X(_02671_));
 sky130_fd_sc_hd__or2_1 _11878_ (.A(_03987_),
    .B(_03998_),
    .X(_02672_));
 sky130_fd_sc_hd__o22ai_4 _11879_ (.A1(_03648_),
    .A2(_03659_),
    .B1(_03670_),
    .B2(_03681_),
    .Y(_02673_));
 sky130_fd_sc_hd__a22oi_4 _11880_ (.A1(net465),
    .A2(net702),
    .B1(net712),
    .B2(net454),
    .Y(_02674_));
 sky130_fd_sc_hd__and4_1 _11881_ (.A(net454),
    .B(net464),
    .C(net702),
    .D(net712),
    .X(_02675_));
 sky130_fd_sc_hd__nor2_2 _11882_ (.A(_02674_),
    .B(_02675_),
    .Y(_02676_));
 sky130_fd_sc_hd__nand2_4 _11883_ (.A(net474),
    .B(net694),
    .Y(_02677_));
 sky130_fd_sc_hd__xnor2_4 _11884_ (.A(_02676_),
    .B(_02677_),
    .Y(_02678_));
 sky130_fd_sc_hd__nand2_2 _11885_ (.A(_02673_),
    .B(_02678_),
    .Y(_02679_));
 sky130_fd_sc_hd__xor2_2 _11886_ (.A(_02673_),
    .B(_02678_),
    .X(_02680_));
 sky130_fd_sc_hd__nand2_2 _11887_ (.A(_02672_),
    .B(_02680_),
    .Y(_02681_));
 sky130_fd_sc_hd__or2_1 _11888_ (.A(_02672_),
    .B(_02680_),
    .X(_02682_));
 sky130_fd_sc_hd__nand2_2 _11889_ (.A(_02681_),
    .B(_02682_),
    .Y(_02683_));
 sky130_fd_sc_hd__o21a_2 _11890_ (.A1(_02670_),
    .A2(_02671_),
    .B1(_02683_),
    .X(_02684_));
 sky130_fd_sc_hd__nor3_4 _11891_ (.A(_02670_),
    .B(_02671_),
    .C(_02683_),
    .Y(_02685_));
 sky130_fd_sc_hd__a211oi_4 _11892_ (.A1(_03888_),
    .A2(_04096_),
    .B1(_02684_),
    .C1(_02685_),
    .Y(_02686_));
 sky130_fd_sc_hd__o211a_1 _11893_ (.A1(_02684_),
    .A2(_02685_),
    .B1(_03888_),
    .C1(_04096_),
    .X(_02687_));
 sky130_fd_sc_hd__a22oi_2 _11894_ (.A1(net518),
    .A2(net651),
    .B1(net659),
    .B2(net509),
    .Y(_02688_));
 sky130_fd_sc_hd__and4_2 _11895_ (.A(net509),
    .B(net517),
    .C(net651),
    .D(net659),
    .X(_02689_));
 sky130_fd_sc_hd__and4bb_2 _11896_ (.A_N(_02688_),
    .B_N(_02689_),
    .C(net526),
    .D(net642),
    .X(_02690_));
 sky130_fd_sc_hd__o2bb2a_1 _11897_ (.A1_N(net526),
    .A2_N(net642),
    .B1(_02688_),
    .B2(_02689_),
    .X(_02691_));
 sky130_fd_sc_hd__nor2_1 _11898_ (.A(_02690_),
    .B(_02691_),
    .Y(_02692_));
 sky130_fd_sc_hd__a22oi_2 _11899_ (.A1(net492),
    .A2(net676),
    .B1(net685),
    .B2(net482),
    .Y(_02693_));
 sky130_fd_sc_hd__and4_1 _11900_ (.A(net482),
    .B(net492),
    .C(net676),
    .D(net685),
    .X(_02694_));
 sky130_fd_sc_hd__nor2_1 _11901_ (.A(_02693_),
    .B(_02694_),
    .Y(_02695_));
 sky130_fd_sc_hd__nand2_2 _11902_ (.A(net502),
    .B(net668),
    .Y(_02696_));
 sky130_fd_sc_hd__xnor2_2 _11903_ (.A(_02695_),
    .B(_02696_),
    .Y(_02697_));
 sky130_fd_sc_hd__o21ba_1 _11904_ (.A1(_04707_),
    .A2(_04740_),
    .B1_N(_04718_),
    .X(_02698_));
 sky130_fd_sc_hd__and2b_2 _11905_ (.A_N(_02698_),
    .B(_02697_),
    .X(_02699_));
 sky130_fd_sc_hd__xnor2_1 _11906_ (.A(_02697_),
    .B(_02698_),
    .Y(_02700_));
 sky130_fd_sc_hd__and2_2 _11907_ (.A(_02692_),
    .B(_02700_),
    .X(_02701_));
 sky130_fd_sc_hd__nor2_1 _11908_ (.A(_02692_),
    .B(_02700_),
    .Y(_02702_));
 sky130_fd_sc_hd__or2_1 _11909_ (.A(_02701_),
    .B(_02702_),
    .X(_02703_));
 sky130_fd_sc_hd__a21o_2 _11910_ (.A1(_04030_),
    .A2(_04052_),
    .B1(_02703_),
    .X(_02704_));
 sky130_fd_sc_hd__nand3_2 _11911_ (.A(_04030_),
    .B(_04052_),
    .C(_02703_),
    .Y(_02705_));
 sky130_fd_sc_hd__o211ai_4 _11912_ (.A1(_04772_),
    .A2(_04794_),
    .B1(_02704_),
    .C1(_02705_),
    .Y(_02706_));
 sky130_fd_sc_hd__a211o_1 _11913_ (.A1(_02704_),
    .A2(_02705_),
    .B1(_04772_),
    .C1(_04794_),
    .X(_02707_));
 sky130_fd_sc_hd__a2bb2o_2 _11914_ (.A1_N(_02686_),
    .A2_N(_02687_),
    .B1(_02706_),
    .B2(_02707_),
    .X(_02708_));
 sky130_fd_sc_hd__or4bb_4 _11915_ (.A(_02686_),
    .B(_02687_),
    .C_N(_02706_),
    .D_N(_02707_),
    .X(_02709_));
 sky130_fd_sc_hd__inv_2 _11916_ (.A(_02709_),
    .Y(_02710_));
 sky130_fd_sc_hd__o211a_4 _11917_ (.A1(_04445_),
    .A2(_04881_),
    .B1(_02708_),
    .C1(_02709_),
    .X(_02711_));
 sky130_fd_sc_hd__a211oi_4 _11918_ (.A1(_02708_),
    .A2(_02709_),
    .B1(_04445_),
    .C1(_04881_),
    .Y(_02712_));
 sky130_fd_sc_hd__a22oi_1 _11919_ (.A1(net326),
    .A2(net870),
    .B1(net880),
    .B2(net317),
    .Y(_02713_));
 sky130_fd_sc_hd__and4_1 _11920_ (.A(net317),
    .B(net326),
    .C(net870),
    .D(net880),
    .X(_02714_));
 sky130_fd_sc_hd__or2_1 _11921_ (.A(_02713_),
    .B(_02714_),
    .X(_02715_));
 sky130_fd_sc_hd__nand2_1 _11922_ (.A(net335),
    .B(net860),
    .Y(_02716_));
 sky130_fd_sc_hd__nor2_2 _11923_ (.A(_02715_),
    .B(_02716_),
    .Y(_02717_));
 sky130_fd_sc_hd__and2_1 _11924_ (.A(_02715_),
    .B(_02716_),
    .X(_02718_));
 sky130_fd_sc_hd__nor2_1 _11925_ (.A(_02717_),
    .B(_02718_),
    .Y(_02719_));
 sky130_fd_sc_hd__a31o_4 _11926_ (.A1(net564),
    .A2(net625),
    .A3(_06246_),
    .B1(_06235_),
    .X(_02720_));
 sky130_fd_sc_hd__a31o_1 _11927_ (.A1(net526),
    .A2(net651),
    .A3(_04674_),
    .B1(_04663_),
    .X(_02721_));
 sky130_fd_sc_hd__nand2_1 _11928_ (.A(net563),
    .B(net625),
    .Y(_02722_));
 sky130_fd_sc_hd__a22oi_2 _11929_ (.A1(net551),
    .A2(net625),
    .B1(net633),
    .B2(net536),
    .Y(_02723_));
 sky130_fd_sc_hd__and4_1 _11930_ (.A(net536),
    .B(net551),
    .C(net625),
    .D(net633),
    .X(_02724_));
 sky130_fd_sc_hd__nor2_2 _11931_ (.A(_02723_),
    .B(_02724_),
    .Y(_02725_));
 sky130_fd_sc_hd__nand2_1 _11932_ (.A(net565),
    .B(net617),
    .Y(_02726_));
 sky130_fd_sc_hd__xnor2_1 _11933_ (.A(_02725_),
    .B(_02726_),
    .Y(_02727_));
 sky130_fd_sc_hd__and2_2 _11934_ (.A(_02721_),
    .B(_02727_),
    .X(_02728_));
 sky130_fd_sc_hd__nor2_1 _11935_ (.A(_02721_),
    .B(_02727_),
    .Y(_02729_));
 sky130_fd_sc_hd__nor2_4 _11936_ (.A(_02728_),
    .B(_02729_),
    .Y(_02730_));
 sky130_fd_sc_hd__xnor2_2 _11937_ (.A(_02720_),
    .B(_02730_),
    .Y(_02731_));
 sky130_fd_sc_hd__a21oi_2 _11938_ (.A1(_06203_),
    .A2(_06290_),
    .B1(_06279_),
    .Y(_02732_));
 sky130_fd_sc_hd__xor2_1 _11939_ (.A(_02731_),
    .B(_02732_),
    .X(_02733_));
 sky130_fd_sc_hd__and2_1 _11940_ (.A(_02719_),
    .B(_02733_),
    .X(_02734_));
 sky130_fd_sc_hd__nor2_1 _11941_ (.A(_02719_),
    .B(_02733_),
    .Y(_02735_));
 sky130_fd_sc_hd__a211o_4 _11942_ (.A1(_04827_),
    .A2(_04849_),
    .B1(_02734_),
    .C1(_02735_),
    .X(_02736_));
 sky130_fd_sc_hd__clkinv_2 _11943_ (.A(_02736_),
    .Y(_02737_));
 sky130_fd_sc_hd__o211a_2 _11944_ (.A1(_02734_),
    .A2(_02735_),
    .B1(_04827_),
    .C1(_04849_),
    .X(_02738_));
 sky130_fd_sc_hd__a211o_4 _11945_ (.A1(_06322_),
    .A2(_06344_),
    .B1(_02737_),
    .C1(_02738_),
    .X(_02739_));
 sky130_fd_sc_hd__o211ai_4 _11946_ (.A1(_02737_),
    .A2(_02738_),
    .B1(_06322_),
    .C1(_06344_),
    .Y(_02740_));
 sky130_fd_sc_hd__and4bb_4 _11947_ (.A_N(_02711_),
    .B_N(_02712_),
    .C(_02739_),
    .D(_02740_),
    .X(_02741_));
 sky130_fd_sc_hd__a2bb2oi_4 _11948_ (.A1_N(_02711_),
    .A2_N(_02712_),
    .B1(_02739_),
    .B2(_02740_),
    .Y(_02742_));
 sky130_fd_sc_hd__a211oi_4 _11949_ (.A1(_05512_),
    .A2(_06431_),
    .B1(_02741_),
    .C1(_02742_),
    .Y(_02743_));
 sky130_fd_sc_hd__o211a_4 _11950_ (.A1(_02741_),
    .A2(_02742_),
    .B1(_05512_),
    .C1(_06431_),
    .X(_02744_));
 sky130_fd_sc_hd__o21ba_2 _11951_ (.A1(_06105_),
    .A2(_06387_),
    .B1_N(_06376_),
    .X(_02745_));
 sky130_fd_sc_hd__a22oi_4 _11952_ (.A1(net372),
    .A2(net810),
    .B1(net821),
    .B2(net363),
    .Y(_02746_));
 sky130_fd_sc_hd__and4_2 _11953_ (.A(net363),
    .B(net372),
    .C(net810),
    .D(net821),
    .X(_02747_));
 sky130_fd_sc_hd__nand2_1 _11954_ (.A(net383),
    .B(net800),
    .Y(_02748_));
 sky130_fd_sc_hd__o21a_1 _11955_ (.A1(_02746_),
    .A2(_02747_),
    .B1(_02748_),
    .X(_02749_));
 sky130_fd_sc_hd__nor3_2 _11956_ (.A(_02746_),
    .B(_02747_),
    .C(_02748_),
    .Y(_02750_));
 sky130_fd_sc_hd__nor2_1 _11957_ (.A(_02749_),
    .B(_02750_),
    .Y(_02751_));
 sky130_fd_sc_hd__or3_1 _11958_ (.A(_08534_),
    .B(_08552_),
    .C(_02751_),
    .X(_02752_));
 sky130_fd_sc_hd__o21ai_1 _11959_ (.A1(_08534_),
    .A2(_08552_),
    .B1(_02751_),
    .Y(_02753_));
 sky130_fd_sc_hd__and2_1 _11960_ (.A(_02752_),
    .B(_02753_),
    .X(_02754_));
 sky130_fd_sc_hd__nand3_1 _11961_ (.A(net388),
    .B(net790),
    .C(_02754_),
    .Y(_02755_));
 sky130_fd_sc_hd__a21o_1 _11962_ (.A1(net388),
    .A2(net790),
    .B1(_02754_),
    .X(_02756_));
 sky130_fd_sc_hd__nand2_1 _11963_ (.A(_02755_),
    .B(_02756_),
    .Y(_02757_));
 sky130_fd_sc_hd__a31o_1 _11964_ (.A1(net388),
    .A2(net800),
    .A3(_08566_),
    .B1(_08565_),
    .X(_02758_));
 sky130_fd_sc_hd__nand2b_2 _11965_ (.A_N(_02757_),
    .B(_02758_),
    .Y(_02759_));
 sky130_fd_sc_hd__nand2b_1 _11966_ (.A_N(_02758_),
    .B(_02757_),
    .Y(_02760_));
 sky130_fd_sc_hd__nand2_1 _11967_ (.A(_02759_),
    .B(_02760_),
    .Y(_02761_));
 sky130_fd_sc_hd__nand2_1 _11968_ (.A(net396),
    .B(net778),
    .Y(_02762_));
 sky130_fd_sc_hd__or2_2 _11969_ (.A(_02761_),
    .B(_02762_),
    .X(_02763_));
 sky130_fd_sc_hd__nand2_1 _11970_ (.A(_02761_),
    .B(_02762_),
    .Y(_02764_));
 sky130_fd_sc_hd__and2_1 _11971_ (.A(_02763_),
    .B(_02764_),
    .X(_02765_));
 sky130_fd_sc_hd__a21o_2 _11972_ (.A1(_08574_),
    .A2(_08582_),
    .B1(_08580_),
    .X(_02766_));
 sky130_fd_sc_hd__a21o_2 _11973_ (.A1(_05867_),
    .A2(_06170_),
    .B1(_05878_),
    .X(_02767_));
 sky130_fd_sc_hd__o21ba_1 _11974_ (.A1(_08575_),
    .A2(_08578_),
    .B1_N(_08576_),
    .X(_02768_));
 sky130_fd_sc_hd__o21ba_2 _11975_ (.A1(_06116_),
    .A2(_06149_),
    .B1_N(_06127_),
    .X(_02769_));
 sky130_fd_sc_hd__a22oi_4 _11976_ (.A1(net349),
    .A2(net840),
    .B1(net850),
    .B2(net340),
    .Y(_02770_));
 sky130_fd_sc_hd__and4_1 _11977_ (.A(net340),
    .B(net349),
    .C(net840),
    .D(net850),
    .X(_02771_));
 sky130_fd_sc_hd__nor2_1 _11978_ (.A(_02770_),
    .B(_02771_),
    .Y(_02772_));
 sky130_fd_sc_hd__nand2_1 _11979_ (.A(net357),
    .B(net830),
    .Y(_02773_));
 sky130_fd_sc_hd__xnor2_1 _11980_ (.A(_02772_),
    .B(_02773_),
    .Y(_02774_));
 sky130_fd_sc_hd__and2b_1 _11981_ (.A_N(_02769_),
    .B(_02774_),
    .X(_02775_));
 sky130_fd_sc_hd__xnor2_1 _11982_ (.A(_02769_),
    .B(_02774_),
    .Y(_02776_));
 sky130_fd_sc_hd__and2b_1 _11983_ (.A_N(_02768_),
    .B(_02776_),
    .X(_02777_));
 sky130_fd_sc_hd__xnor2_1 _11984_ (.A(_02768_),
    .B(_02776_),
    .Y(_02778_));
 sky130_fd_sc_hd__and2b_2 _11985_ (.A_N(_02767_),
    .B(_02778_),
    .X(_02779_));
 sky130_fd_sc_hd__and2b_1 _11986_ (.A_N(_02778_),
    .B(_02767_),
    .X(_02780_));
 sky130_fd_sc_hd__nor2_4 _11987_ (.A(_02779_),
    .B(_02780_),
    .Y(_02781_));
 sky130_fd_sc_hd__xnor2_2 _11988_ (.A(_02766_),
    .B(_02781_),
    .Y(_02782_));
 sky130_fd_sc_hd__a21oi_4 _11989_ (.A1(_08584_),
    .A2(_08587_),
    .B1(_02782_),
    .Y(_02783_));
 sky130_fd_sc_hd__and3_2 _11990_ (.A(_08584_),
    .B(_08587_),
    .C(_02782_),
    .X(_02784_));
 sky130_fd_sc_hd__nor3b_4 _11991_ (.A(_02783_),
    .B(_02784_),
    .C_N(_02765_),
    .Y(_02785_));
 sky130_fd_sc_hd__o21ba_2 _11992_ (.A1(_02783_),
    .A2(_02784_),
    .B1_N(_02765_),
    .X(_02786_));
 sky130_fd_sc_hd__nor3_4 _11993_ (.A(_02745_),
    .B(_02785_),
    .C(_02786_),
    .Y(_02787_));
 sky130_fd_sc_hd__o21a_2 _11994_ (.A1(_02785_),
    .A2(_02786_),
    .B1(_02745_),
    .X(_02788_));
 sky130_fd_sc_hd__a211oi_4 _11995_ (.A1(_08589_),
    .A2(_08591_),
    .B1(_02787_),
    .C1(_02788_),
    .Y(_02789_));
 sky130_fd_sc_hd__o211a_4 _11996_ (.A1(_02787_),
    .A2(_02788_),
    .B1(_08589_),
    .C1(_08591_),
    .X(_02790_));
 sky130_fd_sc_hd__nor4_4 _11997_ (.A(net119),
    .B(_02744_),
    .C(_02789_),
    .D(_02790_),
    .Y(_02791_));
 sky130_fd_sc_hd__or4_4 _11998_ (.A(net119),
    .B(_02744_),
    .C(_02789_),
    .D(_02790_),
    .X(_02792_));
 sky130_fd_sc_hd__o22ai_4 _11999_ (.A1(net119),
    .A2(_02744_),
    .B1(_02789_),
    .B2(_02790_),
    .Y(_02793_));
 sky130_fd_sc_hd__o211a_2 _12000_ (.A1(_07563_),
    .A2(_08598_),
    .B1(_02792_),
    .C1(_02793_),
    .X(_02794_));
 sky130_fd_sc_hd__a211oi_4 _12001_ (.A1(_02792_),
    .A2(_02793_),
    .B1(_07563_),
    .C1(_08598_),
    .Y(_02795_));
 sky130_fd_sc_hd__a211oi_4 _12002_ (.A1(_08593_),
    .A2(_08595_),
    .B1(_02794_),
    .C1(_02795_),
    .Y(_02796_));
 sky130_fd_sc_hd__o211a_1 _12003_ (.A1(_02794_),
    .A2(_02795_),
    .B1(_08593_),
    .C1(_08595_),
    .X(_02797_));
 sky130_fd_sc_hd__nor2_4 _12004_ (.A(_02796_),
    .B(_02797_),
    .Y(_02798_));
 sky130_fd_sc_hd__nand2_2 _12005_ (.A(_00189_),
    .B(_00191_),
    .Y(_02799_));
 sky130_fd_sc_hd__and2_1 _12006_ (.A(_02798_),
    .B(_02799_),
    .X(_02800_));
 sky130_fd_sc_hd__xor2_4 _12007_ (.A(_02798_),
    .B(_02799_),
    .X(_02801_));
 sky130_fd_sc_hd__a31oi_4 _12008_ (.A1(net396),
    .A2(net790),
    .A3(_08571_),
    .B1(_08569_),
    .Y(_02802_));
 sky130_fd_sc_hd__clkinv_4 _12009_ (.A(_02802_),
    .Y(_02803_));
 sky130_fd_sc_hd__xnor2_4 _12010_ (.A(_02801_),
    .B(_02803_),
    .Y(_02804_));
 sky130_fd_sc_hd__a21oi_4 _12011_ (.A1(_00331_),
    .A2(_00332_),
    .B1(_00329_),
    .Y(_02805_));
 sky130_fd_sc_hd__nor2_2 _12012_ (.A(_02804_),
    .B(_02805_),
    .Y(_02806_));
 sky130_fd_sc_hd__and2_1 _12013_ (.A(_02804_),
    .B(_02805_),
    .X(_02807_));
 sky130_fd_sc_hd__nor2_4 _12014_ (.A(_02806_),
    .B(_02807_),
    .Y(_02808_));
 sky130_fd_sc_hd__o21bai_4 _12015_ (.A1(_00472_),
    .A2(_00619_),
    .B1_N(_00473_),
    .Y(_02809_));
 sky130_fd_sc_hd__nand2_2 _12016_ (.A(_00474_),
    .B(_00621_),
    .Y(_02810_));
 sky130_fd_sc_hd__o21ai_4 _12017_ (.A1(_02575_),
    .A2(_02810_),
    .B1(_02809_),
    .Y(_02811_));
 sky130_fd_sc_hd__xnor2_4 _12018_ (.A(_02808_),
    .B(_02811_),
    .Y(_02812_));
 sky130_fd_sc_hd__a21o_1 _12019_ (.A1(net284),
    .A2(net714),
    .B1(_01225_),
    .X(_02813_));
 sky130_fd_sc_hd__nand2_1 _12020_ (.A(net214),
    .B(_02813_),
    .Y(_02814_));
 sky130_fd_sc_hd__and2_1 _12021_ (.A(net284),
    .B(net697),
    .X(_02815_));
 sky130_fd_sc_hd__o21ai_2 _12022_ (.A1(_00974_),
    .A2(_02815_),
    .B1(net214),
    .Y(_02816_));
 sky130_fd_sc_hd__and2_1 _12023_ (.A(net283),
    .B(net679),
    .X(_02817_));
 sky130_fd_sc_hd__o21ai_2 _12024_ (.A1(_00574_),
    .A2(_02817_),
    .B1(net214),
    .Y(_02818_));
 sky130_fd_sc_hd__and2_1 _12025_ (.A(net283),
    .B(net661),
    .X(_02819_));
 sky130_fd_sc_hd__o21ai_2 _12026_ (.A1(_00287_),
    .A2(_02819_),
    .B1(net213),
    .Y(_02820_));
 sky130_fd_sc_hd__mux2_1 _12027_ (.A0(_02818_),
    .A1(_02820_),
    .S(net288),
    .X(_02821_));
 sky130_fd_sc_hd__mux4_2 _12028_ (.A0(_02814_),
    .A1(_02816_),
    .A2(_02818_),
    .A3(_02820_),
    .S0(net290),
    .S1(net297),
    .X(_02822_));
 sky130_fd_sc_hd__nand2_1 _12029_ (.A(_05899_),
    .B(net213),
    .Y(_02823_));
 sky130_fd_sc_hd__a21o_1 _12030_ (.A1(net283),
    .A2(net643),
    .B1(_07987_),
    .X(_02824_));
 sky130_fd_sc_hd__nand2_1 _12031_ (.A(net212),
    .B(_02824_),
    .Y(_02825_));
 sky130_fd_sc_hd__nor2_2 _12032_ (.A(net607),
    .B(_03258_),
    .Y(_02826_));
 sky130_fd_sc_hd__o21ai_1 _12033_ (.A1(_05910_),
    .A2(_02826_),
    .B1(net213),
    .Y(_02827_));
 sky130_fd_sc_hd__mux2_2 _12034_ (.A0(_02825_),
    .A1(_02827_),
    .S(net287),
    .X(_02828_));
 sky130_fd_sc_hd__or3_2 _12035_ (.A(net584),
    .B(net288),
    .C(_02823_),
    .X(_02829_));
 sky130_fd_sc_hd__o21ai_4 _12036_ (.A1(net294),
    .A2(_02828_),
    .B1(_02829_),
    .Y(_02830_));
 sky130_fd_sc_hd__inv_2 _12037_ (.A(_02830_),
    .Y(_02831_));
 sky130_fd_sc_hd__mux2_1 _12038_ (.A0(_02822_),
    .A1(_02831_),
    .S(net300),
    .X(_02832_));
 sky130_fd_sc_hd__mux2_1 _12039_ (.A0(net875),
    .A1(net886),
    .S(net611),
    .X(_02833_));
 sky130_fd_sc_hd__nand2_1 _12040_ (.A(net214),
    .B(_02833_),
    .Y(_02834_));
 sky130_fd_sc_hd__mux2_1 _12041_ (.A0(net855),
    .A1(net868),
    .S(net611),
    .X(_02835_));
 sky130_fd_sc_hd__nand2_1 _12042_ (.A(net214),
    .B(_02835_),
    .Y(_02836_));
 sky130_fd_sc_hd__mux2_1 _12043_ (.A0(net838),
    .A1(net845),
    .S(net611),
    .X(_02837_));
 sky130_fd_sc_hd__nand2_1 _12044_ (.A(net214),
    .B(_02837_),
    .Y(_02838_));
 sky130_fd_sc_hd__a21o_2 _12045_ (.A1(net286),
    .A2(net816),
    .B1(_02072_),
    .X(_02839_));
 sky130_fd_sc_hd__nand2_1 _12046_ (.A(net215),
    .B(_02839_),
    .Y(_02840_));
 sky130_fd_sc_hd__mux4_2 _12047_ (.A0(_02834_),
    .A1(_02836_),
    .A2(_02838_),
    .A3(_02840_),
    .S0(net291),
    .S1(net296),
    .X(_02841_));
 sky130_fd_sc_hd__mux2_1 _12048_ (.A0(net796),
    .A1(net807),
    .S(net608),
    .X(_02842_));
 sky130_fd_sc_hd__nand2_1 _12049_ (.A(net215),
    .B(_02842_),
    .Y(_02843_));
 sky130_fd_sc_hd__mux2_1 _12050_ (.A0(net771),
    .A1(net780),
    .S(net608),
    .X(_02844_));
 sky130_fd_sc_hd__nand2_1 _12051_ (.A(net215),
    .B(_02844_),
    .Y(_02845_));
 sky130_fd_sc_hd__a21o_1 _12052_ (.A1(net283),
    .A2(net750),
    .B1(_01580_),
    .X(_02846_));
 sky130_fd_sc_hd__nand2_1 _12053_ (.A(net214),
    .B(_02846_),
    .Y(_02847_));
 sky130_fd_sc_hd__and2_2 _12054_ (.A(net284),
    .B(net732),
    .X(_02848_));
 sky130_fd_sc_hd__o21ai_4 _12055_ (.A1(_01451_),
    .A2(_02848_),
    .B1(net214),
    .Y(_02849_));
 sky130_fd_sc_hd__mux4_1 _12056_ (.A0(_02843_),
    .A1(_02845_),
    .A2(_02847_),
    .A3(_02849_),
    .S0(net291),
    .S1(net296),
    .X(_02850_));
 sky130_fd_sc_hd__mux2_1 _12057_ (.A0(_02841_),
    .A1(_02850_),
    .S(net301),
    .X(_02851_));
 sky130_fd_sc_hd__mux2_1 _12058_ (.A0(_02832_),
    .A1(_02851_),
    .S(net552),
    .X(_02852_));
 sky130_fd_sc_hd__or3b_2 _12059_ (.A(net611),
    .B(_03302_),
    .C_N(net215),
    .X(_02853_));
 sky130_fd_sc_hd__mux2_1 _12060_ (.A0(net900),
    .A1(net902),
    .S(net611),
    .X(_02854_));
 sky130_fd_sc_hd__nand2_1 _12061_ (.A(net214),
    .B(_02854_),
    .Y(_02855_));
 sky130_fd_sc_hd__mux2_1 _12062_ (.A0(_02853_),
    .A1(_02855_),
    .S(net291),
    .X(_02856_));
 sky130_fd_sc_hd__or3_4 _12063_ (.A(net577),
    .B(net585),
    .C(_02856_),
    .X(_02857_));
 sky130_fd_sc_hd__o21a_1 _12064_ (.A1(net552),
    .A2(_02857_),
    .B1(net540),
    .X(_02858_));
 sky130_fd_sc_hd__a211o_1 _12065_ (.A1(_03193_),
    .A2(_02852_),
    .B1(_02858_),
    .C1(_02642_),
    .X(_02859_));
 sky130_fd_sc_hd__o21ai_1 _12066_ (.A1(net255),
    .A2(_02812_),
    .B1(_02859_),
    .Y(_08664_));
 sky130_fd_sc_hd__a22o_1 _12067_ (.A1(net420),
    .A2(net738),
    .B1(net756),
    .B2(net404),
    .X(_02860_));
 sky130_fd_sc_hd__and4_1 _12068_ (.A(net404),
    .B(net420),
    .C(net738),
    .D(net756),
    .X(_02861_));
 sky130_fd_sc_hd__inv_2 _12069_ (.A(_02861_),
    .Y(_02862_));
 sky130_fd_sc_hd__and4_1 _12070_ (.A(net413),
    .B(net747),
    .C(_02860_),
    .D(_02862_),
    .X(_02863_));
 sky130_fd_sc_hd__a22oi_1 _12071_ (.A1(net413),
    .A2(net747),
    .B1(_02860_),
    .B2(_02862_),
    .Y(_02864_));
 sky130_fd_sc_hd__nor2_1 _12072_ (.A(_02863_),
    .B(_02864_),
    .Y(_02865_));
 sky130_fd_sc_hd__o21ba_1 _12073_ (.A1(_02652_),
    .A2(_02655_),
    .B1_N(_02653_),
    .X(_02866_));
 sky130_fd_sc_hd__and2b_2 _12074_ (.A_N(_02866_),
    .B(_02865_),
    .X(_02867_));
 sky130_fd_sc_hd__xnor2_1 _12075_ (.A(_02865_),
    .B(_02866_),
    .Y(_02868_));
 sky130_fd_sc_hd__a22oi_4 _12076_ (.A1(net436),
    .A2(net721),
    .B1(net730),
    .B2(net428),
    .Y(_02869_));
 sky130_fd_sc_hd__and4_1 _12077_ (.A(net428),
    .B(net436),
    .C(net721),
    .D(net730),
    .X(_02870_));
 sky130_fd_sc_hd__nor2_1 _12078_ (.A(_02869_),
    .B(_02870_),
    .Y(_02871_));
 sky130_fd_sc_hd__nand2_1 _12079_ (.A(net446),
    .B(net712),
    .Y(_02872_));
 sky130_fd_sc_hd__xnor2_1 _12080_ (.A(_02871_),
    .B(_02872_),
    .Y(_02873_));
 sky130_fd_sc_hd__and2_2 _12081_ (.A(_02868_),
    .B(_02873_),
    .X(_02874_));
 sky130_fd_sc_hd__nor2_1 _12082_ (.A(_02868_),
    .B(_02873_),
    .Y(_02875_));
 sky130_fd_sc_hd__or2_2 _12083_ (.A(_02874_),
    .B(_02875_),
    .X(_02876_));
 sky130_fd_sc_hd__a21o_4 _12084_ (.A1(_02658_),
    .A2(_02667_),
    .B1(_02876_),
    .X(_02877_));
 sky130_fd_sc_hd__nand3_4 _12085_ (.A(_02658_),
    .B(_02667_),
    .C(_02876_),
    .Y(_02878_));
 sky130_fd_sc_hd__o21ba_4 _12086_ (.A1(_02674_),
    .A2(_02677_),
    .B1_N(_02675_),
    .X(_02879_));
 sky130_fd_sc_hd__a22oi_4 _12087_ (.A1(net464),
    .A2(net695),
    .B1(net703),
    .B2(net454),
    .Y(_02880_));
 sky130_fd_sc_hd__and4_1 _12088_ (.A(net454),
    .B(net464),
    .C(net695),
    .D(net703),
    .X(_02881_));
 sky130_fd_sc_hd__nor2_1 _12089_ (.A(_02880_),
    .B(_02881_),
    .Y(_02882_));
 sky130_fd_sc_hd__nand2_2 _12090_ (.A(net474),
    .B(net686),
    .Y(_02883_));
 sky130_fd_sc_hd__xnor2_2 _12091_ (.A(_02882_),
    .B(_02883_),
    .Y(_02884_));
 sky130_fd_sc_hd__o21ai_4 _12092_ (.A1(_02661_),
    .A2(_02664_),
    .B1(_02884_),
    .Y(_02885_));
 sky130_fd_sc_hd__or3_1 _12093_ (.A(_02661_),
    .B(_02664_),
    .C(_02884_),
    .X(_02886_));
 sky130_fd_sc_hd__and2_2 _12094_ (.A(_02885_),
    .B(_02886_),
    .X(_02887_));
 sky130_fd_sc_hd__nand2b_2 _12095_ (.A_N(_02879_),
    .B(_02887_),
    .Y(_02888_));
 sky130_fd_sc_hd__xnor2_4 _12096_ (.A(_02879_),
    .B(_02887_),
    .Y(_02889_));
 sky130_fd_sc_hd__a21o_2 _12097_ (.A1(_02877_),
    .A2(_02878_),
    .B1(_02889_),
    .X(_02890_));
 sky130_fd_sc_hd__nand3_4 _12098_ (.A(_02877_),
    .B(_02878_),
    .C(_02889_),
    .Y(_02891_));
 sky130_fd_sc_hd__o211ai_4 _12099_ (.A1(_02670_),
    .A2(_02685_),
    .B1(_02890_),
    .C1(_02891_),
    .Y(_02892_));
 sky130_fd_sc_hd__a211o_2 _12100_ (.A1(_02890_),
    .A2(_02891_),
    .B1(_02670_),
    .C1(_02685_),
    .X(_02893_));
 sky130_fd_sc_hd__a22oi_1 _12101_ (.A1(net519),
    .A2(net643),
    .B1(net652),
    .B2(net509),
    .Y(_02894_));
 sky130_fd_sc_hd__and4_1 _12102_ (.A(net509),
    .B(net519),
    .C(net643),
    .D(net652),
    .X(_02895_));
 sky130_fd_sc_hd__nor2_1 _12103_ (.A(_02894_),
    .B(_02895_),
    .Y(_02896_));
 sky130_fd_sc_hd__nand2_1 _12104_ (.A(net525),
    .B(net633),
    .Y(_02897_));
 sky130_fd_sc_hd__xnor2_1 _12105_ (.A(_02896_),
    .B(_02897_),
    .Y(_02898_));
 sky130_fd_sc_hd__a22oi_2 _12106_ (.A1(net494),
    .A2(net668),
    .B1(net678),
    .B2(net484),
    .Y(_02899_));
 sky130_fd_sc_hd__and4_1 _12107_ (.A(net484),
    .B(net494),
    .C(net668),
    .D(net678),
    .X(_02900_));
 sky130_fd_sc_hd__nor2_1 _12108_ (.A(_02899_),
    .B(_02900_),
    .Y(_02901_));
 sky130_fd_sc_hd__nand2_2 _12109_ (.A(net503),
    .B(net660),
    .Y(_02902_));
 sky130_fd_sc_hd__xnor2_2 _12110_ (.A(_02901_),
    .B(_02902_),
    .Y(_02903_));
 sky130_fd_sc_hd__o21ba_1 _12111_ (.A1(_02693_),
    .A2(_02696_),
    .B1_N(_02694_),
    .X(_02904_));
 sky130_fd_sc_hd__and2b_2 _12112_ (.A_N(_02904_),
    .B(_02903_),
    .X(_02905_));
 sky130_fd_sc_hd__xnor2_1 _12113_ (.A(_02903_),
    .B(_02904_),
    .Y(_02906_));
 sky130_fd_sc_hd__and2_2 _12114_ (.A(_02898_),
    .B(_02906_),
    .X(_02907_));
 sky130_fd_sc_hd__nor2_1 _12115_ (.A(_02898_),
    .B(_02906_),
    .Y(_02908_));
 sky130_fd_sc_hd__or2_2 _12116_ (.A(_02907_),
    .B(_02908_),
    .X(_02909_));
 sky130_fd_sc_hd__a21o_4 _12117_ (.A1(_02679_),
    .A2(_02681_),
    .B1(_02909_),
    .X(_02910_));
 sky130_fd_sc_hd__nand3_2 _12118_ (.A(_02679_),
    .B(_02681_),
    .C(_02909_),
    .Y(_02911_));
 sky130_fd_sc_hd__o211ai_4 _12119_ (.A1(_02699_),
    .A2(_02701_),
    .B1(_02910_),
    .C1(_02911_),
    .Y(_02912_));
 sky130_fd_sc_hd__a211o_2 _12120_ (.A1(_02910_),
    .A2(_02911_),
    .B1(_02699_),
    .C1(_02701_),
    .X(_02913_));
 sky130_fd_sc_hd__a22o_2 _12121_ (.A1(_02892_),
    .A2(_02893_),
    .B1(_02912_),
    .B2(_02913_),
    .X(_02914_));
 sky130_fd_sc_hd__nand4_4 _12122_ (.A(_02892_),
    .B(_02893_),
    .C(_02912_),
    .D(_02913_),
    .Y(_02915_));
 sky130_fd_sc_hd__o211ai_4 _12123_ (.A1(_02686_),
    .A2(_02710_),
    .B1(_02914_),
    .C1(_02915_),
    .Y(_02916_));
 sky130_fd_sc_hd__a211o_2 _12124_ (.A1(_02914_),
    .A2(_02915_),
    .B1(_02686_),
    .C1(_02710_),
    .X(_02917_));
 sky130_fd_sc_hd__o21ba_4 _12125_ (.A1(_02731_),
    .A2(_02732_),
    .B1_N(_02734_),
    .X(_02918_));
 sky130_fd_sc_hd__a22oi_1 _12126_ (.A1(net327),
    .A2(net860),
    .B1(net870),
    .B2(net317),
    .Y(_02919_));
 sky130_fd_sc_hd__and4_1 _12127_ (.A(net317),
    .B(net327),
    .C(net860),
    .D(net871),
    .X(_02920_));
 sky130_fd_sc_hd__or2_1 _12128_ (.A(_02919_),
    .B(_02920_),
    .X(_02921_));
 sky130_fd_sc_hd__nand2_1 _12129_ (.A(net335),
    .B(net850),
    .Y(_02922_));
 sky130_fd_sc_hd__nor2_1 _12130_ (.A(_02921_),
    .B(_02922_),
    .Y(_02923_));
 sky130_fd_sc_hd__and2_1 _12131_ (.A(_02921_),
    .B(_02922_),
    .X(_02924_));
 sky130_fd_sc_hd__nor2_1 _12132_ (.A(_02923_),
    .B(_02924_),
    .Y(_02925_));
 sky130_fd_sc_hd__a31o_4 _12133_ (.A1(net565),
    .A2(net617),
    .A3(_02725_),
    .B1(_02724_),
    .X(_02926_));
 sky130_fd_sc_hd__o2bb2a_1 _12134_ (.A1_N(net554),
    .A2_N(net618),
    .B1(_03258_),
    .B2(_03193_),
    .X(_02927_));
 sky130_fd_sc_hd__and4_1 _12135_ (.A(net540),
    .B(net554),
    .C(net618),
    .D(net625),
    .X(_02928_));
 sky130_fd_sc_hd__nor2_2 _12136_ (.A(_02927_),
    .B(_02928_),
    .Y(_02929_));
 sky130_fd_sc_hd__o21ai_2 _12137_ (.A1(_02689_),
    .A2(_02690_),
    .B1(_02929_),
    .Y(_02930_));
 sky130_fd_sc_hd__or3_1 _12138_ (.A(_02689_),
    .B(_02690_),
    .C(_02929_),
    .X(_02931_));
 sky130_fd_sc_hd__and2_2 _12139_ (.A(_02930_),
    .B(_02931_),
    .X(_02932_));
 sky130_fd_sc_hd__nand2_1 _12140_ (.A(_02926_),
    .B(_02932_),
    .Y(_02933_));
 sky130_fd_sc_hd__xnor2_4 _12141_ (.A(_02926_),
    .B(_02932_),
    .Y(_02934_));
 sky130_fd_sc_hd__a21oi_4 _12142_ (.A1(_02720_),
    .A2(_02730_),
    .B1(_02728_),
    .Y(_02935_));
 sky130_fd_sc_hd__xor2_2 _12143_ (.A(_02934_),
    .B(_02935_),
    .X(_02936_));
 sky130_fd_sc_hd__nand2_2 _12144_ (.A(_02925_),
    .B(_02936_),
    .Y(_02937_));
 sky130_fd_sc_hd__or2_1 _12145_ (.A(_02925_),
    .B(_02936_),
    .X(_02938_));
 sky130_fd_sc_hd__nand2_1 _12146_ (.A(_02937_),
    .B(_02938_),
    .Y(_02939_));
 sky130_fd_sc_hd__a21oi_2 _12147_ (.A1(_02704_),
    .A2(_02706_),
    .B1(_02939_),
    .Y(_02940_));
 sky130_fd_sc_hd__and3_1 _12148_ (.A(_02704_),
    .B(_02706_),
    .C(_02939_),
    .X(_02941_));
 sky130_fd_sc_hd__nor2_2 _12149_ (.A(_02940_),
    .B(_02941_),
    .Y(_02942_));
 sky130_fd_sc_hd__xnor2_4 _12150_ (.A(_02918_),
    .B(_02942_),
    .Y(_02943_));
 sky130_fd_sc_hd__nand3_4 _12151_ (.A(_02916_),
    .B(_02917_),
    .C(_02943_),
    .Y(_02944_));
 sky130_fd_sc_hd__a21o_2 _12152_ (.A1(_02916_),
    .A2(_02917_),
    .B1(_02943_),
    .X(_02945_));
 sky130_fd_sc_hd__o211ai_4 _12153_ (.A1(_02711_),
    .A2(_02741_),
    .B1(_02944_),
    .C1(_02945_),
    .Y(_02946_));
 sky130_fd_sc_hd__a211o_2 _12154_ (.A1(_02944_),
    .A2(_02945_),
    .B1(_02711_),
    .C1(_02741_),
    .X(_02947_));
 sky130_fd_sc_hd__nor2_4 _12155_ (.A(_02783_),
    .B(_02785_),
    .Y(_02948_));
 sky130_fd_sc_hd__nand2_4 _12156_ (.A(_02736_),
    .B(_02739_),
    .Y(_02949_));
 sky130_fd_sc_hd__a22oi_4 _12157_ (.A1(net373),
    .A2(net800),
    .B1(net810),
    .B2(net364),
    .Y(_02950_));
 sky130_fd_sc_hd__and4_2 _12158_ (.A(net364),
    .B(net373),
    .C(net800),
    .D(net810),
    .X(_02951_));
 sky130_fd_sc_hd__nand2_1 _12159_ (.A(net383),
    .B(net789),
    .Y(_02952_));
 sky130_fd_sc_hd__o21a_1 _12160_ (.A1(_02950_),
    .A2(_02951_),
    .B1(_02952_),
    .X(_02953_));
 sky130_fd_sc_hd__nor3_2 _12161_ (.A(_02950_),
    .B(_02951_),
    .C(_02952_),
    .Y(_02954_));
 sky130_fd_sc_hd__nor2_1 _12162_ (.A(_02953_),
    .B(_02954_),
    .Y(_02955_));
 sky130_fd_sc_hd__nor3_1 _12163_ (.A(_02747_),
    .B(_02750_),
    .C(_02955_),
    .Y(_02956_));
 sky130_fd_sc_hd__o21a_1 _12164_ (.A1(_02747_),
    .A2(_02750_),
    .B1(_02955_),
    .X(_02957_));
 sky130_fd_sc_hd__nor2_1 _12165_ (.A(_02956_),
    .B(_02957_),
    .Y(_02958_));
 sky130_fd_sc_hd__nand2_1 _12166_ (.A(net388),
    .B(net778),
    .Y(_02959_));
 sky130_fd_sc_hd__xor2_1 _12167_ (.A(_02958_),
    .B(_02959_),
    .X(_02960_));
 sky130_fd_sc_hd__a21oi_1 _12168_ (.A1(_02753_),
    .A2(_02755_),
    .B1(_02960_),
    .Y(_02961_));
 sky130_fd_sc_hd__and3_1 _12169_ (.A(_02753_),
    .B(_02755_),
    .C(_02960_),
    .X(_02962_));
 sky130_fd_sc_hd__nor2_1 _12170_ (.A(_02961_),
    .B(_02962_),
    .Y(_02963_));
 sky130_fd_sc_hd__nand2_1 _12171_ (.A(net396),
    .B(net766),
    .Y(_02964_));
 sky130_fd_sc_hd__xnor2_1 _12172_ (.A(_02963_),
    .B(_02964_),
    .Y(_02965_));
 sky130_fd_sc_hd__a22oi_2 _12173_ (.A1(net349),
    .A2(net830),
    .B1(net840),
    .B2(net341),
    .Y(_02966_));
 sky130_fd_sc_hd__and4_1 _12174_ (.A(net341),
    .B(net349),
    .C(net830),
    .D(net840),
    .X(_02967_));
 sky130_fd_sc_hd__nor2_1 _12175_ (.A(_02966_),
    .B(_02967_),
    .Y(_02968_));
 sky130_fd_sc_hd__nand2_2 _12176_ (.A(net357),
    .B(net821),
    .Y(_02969_));
 sky130_fd_sc_hd__xnor2_2 _12177_ (.A(_02968_),
    .B(_02969_),
    .Y(_02970_));
 sky130_fd_sc_hd__o21a_1 _12178_ (.A1(_02714_),
    .A2(_02717_),
    .B1(_02970_),
    .X(_02971_));
 sky130_fd_sc_hd__nor3_2 _12179_ (.A(_02714_),
    .B(_02717_),
    .C(_02970_),
    .Y(_02972_));
 sky130_fd_sc_hd__nor2_4 _12180_ (.A(_02971_),
    .B(_02972_),
    .Y(_02973_));
 sky130_fd_sc_hd__o21ba_4 _12181_ (.A1(_02770_),
    .A2(_02773_),
    .B1_N(_02771_),
    .X(_02974_));
 sky130_fd_sc_hd__xor2_4 _12182_ (.A(_02973_),
    .B(_02974_),
    .X(_02975_));
 sky130_fd_sc_hd__nor2_4 _12183_ (.A(_02775_),
    .B(_02777_),
    .Y(_02976_));
 sky130_fd_sc_hd__xnor2_4 _12184_ (.A(_02975_),
    .B(_02976_),
    .Y(_02977_));
 sky130_fd_sc_hd__a21oi_4 _12185_ (.A1(_02766_),
    .A2(_02781_),
    .B1(_02779_),
    .Y(_02978_));
 sky130_fd_sc_hd__xor2_2 _12186_ (.A(_02977_),
    .B(_02978_),
    .X(_02979_));
 sky130_fd_sc_hd__nand2_2 _12187_ (.A(_02965_),
    .B(_02979_),
    .Y(_02980_));
 sky130_fd_sc_hd__or2_1 _12188_ (.A(_02965_),
    .B(_02979_),
    .X(_02981_));
 sky130_fd_sc_hd__nand2_2 _12189_ (.A(_02980_),
    .B(_02981_),
    .Y(_02982_));
 sky130_fd_sc_hd__xnor2_4 _12190_ (.A(_02949_),
    .B(_02982_),
    .Y(_02983_));
 sky130_fd_sc_hd__and2b_1 _12191_ (.A_N(_02948_),
    .B(_02983_),
    .X(_02984_));
 sky130_fd_sc_hd__xnor2_4 _12192_ (.A(_02948_),
    .B(_02983_),
    .Y(_02985_));
 sky130_fd_sc_hd__nand3_4 _12193_ (.A(_02946_),
    .B(_02947_),
    .C(_02985_),
    .Y(_02986_));
 sky130_fd_sc_hd__a21o_2 _12194_ (.A1(_02946_),
    .A2(_02947_),
    .B1(_02985_),
    .X(_02987_));
 sky130_fd_sc_hd__o211a_2 _12195_ (.A1(_02743_),
    .A2(_02791_),
    .B1(_02986_),
    .C1(_02987_),
    .X(_02988_));
 sky130_fd_sc_hd__a211oi_4 _12196_ (.A1(_02986_),
    .A2(_02987_),
    .B1(_02743_),
    .C1(_02791_),
    .Y(_02989_));
 sky130_fd_sc_hd__nor2_2 _12197_ (.A(_02787_),
    .B(_02789_),
    .Y(_02990_));
 sky130_fd_sc_hd__or3_4 _12198_ (.A(_02988_),
    .B(_02989_),
    .C(_02990_),
    .X(_02991_));
 sky130_fd_sc_hd__o21ai_4 _12199_ (.A1(_02988_),
    .A2(_02989_),
    .B1(_02990_),
    .Y(_02992_));
 sky130_fd_sc_hd__or2_2 _12200_ (.A(_02794_),
    .B(_02796_),
    .X(_02993_));
 sky130_fd_sc_hd__and3_4 _12201_ (.A(_02991_),
    .B(_02992_),
    .C(_02993_),
    .X(_02994_));
 sky130_fd_sc_hd__a21oi_4 _12202_ (.A1(_02991_),
    .A2(_02992_),
    .B1(_02993_),
    .Y(_02995_));
 sky130_fd_sc_hd__a211oi_4 _12203_ (.A1(_02759_),
    .A2(_02763_),
    .B1(_02994_),
    .C1(_02995_),
    .Y(_02996_));
 sky130_fd_sc_hd__o211a_2 _12204_ (.A1(_02994_),
    .A2(_02995_),
    .B1(_02759_),
    .C1(_02763_),
    .X(_02997_));
 sky130_fd_sc_hd__a21oi_4 _12205_ (.A1(_02801_),
    .A2(_02803_),
    .B1(_02800_),
    .Y(_02998_));
 sky130_fd_sc_hd__nor3_4 _12206_ (.A(_02996_),
    .B(_02997_),
    .C(_02998_),
    .Y(_02999_));
 sky130_fd_sc_hd__o21a_4 _12207_ (.A1(_02996_),
    .A2(_02997_),
    .B1(_02998_),
    .X(_03000_));
 sky130_fd_sc_hd__nor2_2 _12208_ (.A(_02999_),
    .B(_03000_),
    .Y(_03001_));
 sky130_fd_sc_hd__a21o_1 _12209_ (.A1(_02808_),
    .A2(_02811_),
    .B1(_02806_),
    .X(_03002_));
 sky130_fd_sc_hd__xnor2_2 _12210_ (.A(_03001_),
    .B(_03002_),
    .Y(_03003_));
 sky130_fd_sc_hd__mux2_1 _12211_ (.A0(_02599_),
    .A1(_02602_),
    .S(net287),
    .X(_03004_));
 sky130_fd_sc_hd__mux2_1 _12212_ (.A0(_02604_),
    .A1(_02609_),
    .S(net288),
    .X(_03005_));
 sky130_fd_sc_hd__mux2_1 _12213_ (.A0(_03004_),
    .A1(_03005_),
    .S(net294),
    .X(_03006_));
 sky130_fd_sc_hd__nor2_1 _12214_ (.A(net598),
    .B(_02607_),
    .Y(_03007_));
 sky130_fd_sc_hd__a21oi_1 _12215_ (.A1(net598),
    .A2(_02611_),
    .B1(_03007_),
    .Y(_03008_));
 sky130_fd_sc_hd__inv_2 _12216_ (.A(_03008_),
    .Y(_03009_));
 sky130_fd_sc_hd__nor2_4 _12217_ (.A(net293),
    .B(_03009_),
    .Y(_03010_));
 sky130_fd_sc_hd__inv_2 _12218_ (.A(_03010_),
    .Y(_03011_));
 sky130_fd_sc_hd__mux2_1 _12219_ (.A0(_03006_),
    .A1(_03011_),
    .S(net300),
    .X(_03012_));
 sky130_fd_sc_hd__mux2_1 _12220_ (.A0(_02621_),
    .A1(_02624_),
    .S(net288),
    .X(_03013_));
 sky130_fd_sc_hd__mux2_1 _12221_ (.A0(_02626_),
    .A1(_02630_),
    .S(net287),
    .X(_03014_));
 sky130_fd_sc_hd__mux2_1 _12222_ (.A0(_03013_),
    .A1(_03014_),
    .S(net293),
    .X(_03015_));
 sky130_fd_sc_hd__mux2_1 _12223_ (.A0(_02632_),
    .A1(_02635_),
    .S(net288),
    .X(_03016_));
 sky130_fd_sc_hd__mux2_1 _12224_ (.A0(_02597_),
    .A1(_02637_),
    .S(net596),
    .X(_03017_));
 sky130_fd_sc_hd__mux2_1 _12225_ (.A0(_03016_),
    .A1(_03017_),
    .S(net294),
    .X(_03018_));
 sky130_fd_sc_hd__mux2_1 _12226_ (.A0(_03015_),
    .A1(_03018_),
    .S(net300),
    .X(_03019_));
 sky130_fd_sc_hd__mux2_1 _12227_ (.A0(_03012_),
    .A1(_03019_),
    .S(net554),
    .X(_03020_));
 sky130_fd_sc_hd__mux2_2 _12228_ (.A0(_02619_),
    .A1(_02646_),
    .S(net597),
    .X(_03021_));
 sky130_fd_sc_hd__or3_4 _12229_ (.A(net566),
    .B(net584),
    .C(_03021_),
    .X(_03022_));
 sky130_fd_sc_hd__or2_1 _12230_ (.A(net206),
    .B(_03022_),
    .X(_03023_));
 sky130_fd_sc_hd__a22o_1 _12231_ (.A1(_03193_),
    .A2(_03020_),
    .B1(_03023_),
    .B2(net209),
    .X(_03024_));
 sky130_fd_sc_hd__o21ai_1 _12232_ (.A1(net255),
    .A2(_03003_),
    .B1(_03024_),
    .Y(_08675_));
 sky130_fd_sc_hd__and2_4 _12233_ (.A(net426),
    .B(net736),
    .X(_03025_));
 sky130_fd_sc_hd__a21oi_4 _12234_ (.A1(net410),
    .A2(net751),
    .B1(_03025_),
    .Y(_03026_));
 sky130_fd_sc_hd__and3_4 _12235_ (.A(net410),
    .B(net751),
    .C(_03025_),
    .X(_03027_));
 sky130_fd_sc_hd__nor2_8 _12236_ (.A(_03026_),
    .B(_03027_),
    .Y(_03028_));
 sky130_fd_sc_hd__nand2_2 _12237_ (.A(net413),
    .B(net738),
    .Y(_03029_));
 sky130_fd_sc_hd__xnor2_4 _12238_ (.A(_03028_),
    .B(_03029_),
    .Y(_03030_));
 sky130_fd_sc_hd__nor2_2 _12239_ (.A(_02861_),
    .B(_02863_),
    .Y(_03031_));
 sky130_fd_sc_hd__nand2b_2 _12240_ (.A_N(_03031_),
    .B(_03030_),
    .Y(_03032_));
 sky130_fd_sc_hd__xor2_4 _12241_ (.A(_03030_),
    .B(_03031_),
    .X(_03033_));
 sky130_fd_sc_hd__a22oi_1 _12242_ (.A1(net436),
    .A2(net712),
    .B1(net721),
    .B2(net428),
    .Y(_03034_));
 sky130_fd_sc_hd__and4_2 _12243_ (.A(net428),
    .B(net436),
    .C(net712),
    .D(net721),
    .X(_03035_));
 sky130_fd_sc_hd__or2_1 _12244_ (.A(_03034_),
    .B(_03035_),
    .X(_03036_));
 sky130_fd_sc_hd__nand2_1 _12245_ (.A(net446),
    .B(net703),
    .Y(_03037_));
 sky130_fd_sc_hd__nor2_2 _12246_ (.A(_03036_),
    .B(_03037_),
    .Y(_03038_));
 sky130_fd_sc_hd__nand2_1 _12247_ (.A(_03036_),
    .B(_03037_),
    .Y(_03039_));
 sky130_fd_sc_hd__and2b_4 _12248_ (.A_N(_03038_),
    .B(_03039_),
    .X(_03040_));
 sky130_fd_sc_hd__nand2b_2 _12249_ (.A_N(_03033_),
    .B(_03040_),
    .Y(_03041_));
 sky130_fd_sc_hd__xnor2_4 _12250_ (.A(_03033_),
    .B(_03040_),
    .Y(_03042_));
 sky130_fd_sc_hd__o21ai_4 _12251_ (.A1(_02867_),
    .A2(_02874_),
    .B1(_03042_),
    .Y(_03043_));
 sky130_fd_sc_hd__or3_4 _12252_ (.A(_02867_),
    .B(_02874_),
    .C(_03042_),
    .X(_03044_));
 sky130_fd_sc_hd__o21ba_4 _12253_ (.A1(_02880_),
    .A2(_02883_),
    .B1_N(_02881_),
    .X(_03045_));
 sky130_fd_sc_hd__o21ba_4 _12254_ (.A1(_02869_),
    .A2(_02872_),
    .B1_N(_02870_),
    .X(_03046_));
 sky130_fd_sc_hd__a22oi_4 _12255_ (.A1(net472),
    .A2(net686),
    .B1(net695),
    .B2(net455),
    .Y(_03047_));
 sky130_fd_sc_hd__and4_1 _12256_ (.A(net455),
    .B(net472),
    .C(net686),
    .D(net695),
    .X(_03048_));
 sky130_fd_sc_hd__nor2_2 _12257_ (.A(_03047_),
    .B(_03048_),
    .Y(_03049_));
 sky130_fd_sc_hd__nand2_4 _12258_ (.A(net479),
    .B(net678),
    .Y(_03050_));
 sky130_fd_sc_hd__xnor2_4 _12259_ (.A(_03049_),
    .B(_03050_),
    .Y(_03051_));
 sky130_fd_sc_hd__nand2b_1 _12260_ (.A_N(_03046_),
    .B(_03051_),
    .Y(_03052_));
 sky130_fd_sc_hd__xnor2_4 _12261_ (.A(_03046_),
    .B(_03051_),
    .Y(_03053_));
 sky130_fd_sc_hd__nand2b_1 _12262_ (.A_N(_03045_),
    .B(_03053_),
    .Y(_03054_));
 sky130_fd_sc_hd__xnor2_4 _12263_ (.A(_03045_),
    .B(_03053_),
    .Y(_03055_));
 sky130_fd_sc_hd__a21o_1 _12264_ (.A1(_03043_),
    .A2(_03044_),
    .B1(_03055_),
    .X(_03056_));
 sky130_fd_sc_hd__nand3_4 _12265_ (.A(_03043_),
    .B(_03044_),
    .C(_03055_),
    .Y(_03057_));
 sky130_fd_sc_hd__nand2_2 _12266_ (.A(_03056_),
    .B(_03057_),
    .Y(_03058_));
 sky130_fd_sc_hd__a21oi_4 _12267_ (.A1(_02877_),
    .A2(_02891_),
    .B1(_03058_),
    .Y(_03059_));
 sky130_fd_sc_hd__and3_2 _12268_ (.A(_02877_),
    .B(_02891_),
    .C(_03058_),
    .X(_03060_));
 sky130_fd_sc_hd__a22oi_4 _12269_ (.A1(net519),
    .A2(net634),
    .B1(net642),
    .B2(net511),
    .Y(_03061_));
 sky130_fd_sc_hd__and4_1 _12270_ (.A(net511),
    .B(net519),
    .C(net634),
    .D(net643),
    .X(_03062_));
 sky130_fd_sc_hd__nor2_1 _12271_ (.A(_03061_),
    .B(_03062_),
    .Y(_03063_));
 sky130_fd_sc_hd__nand2_1 _12272_ (.A(net528),
    .B(net625),
    .Y(_03064_));
 sky130_fd_sc_hd__xnor2_1 _12273_ (.A(_03063_),
    .B(_03064_),
    .Y(_03065_));
 sky130_fd_sc_hd__a22oi_2 _12274_ (.A1(net494),
    .A2(net660),
    .B1(net668),
    .B2(net484),
    .Y(_03066_));
 sky130_fd_sc_hd__and4_1 _12275_ (.A(net484),
    .B(net494),
    .C(net660),
    .D(net668),
    .X(_03067_));
 sky130_fd_sc_hd__nor2_1 _12276_ (.A(_03066_),
    .B(_03067_),
    .Y(_03068_));
 sky130_fd_sc_hd__nand2_2 _12277_ (.A(net503),
    .B(net652),
    .Y(_03069_));
 sky130_fd_sc_hd__xnor2_2 _12278_ (.A(_03068_),
    .B(_03069_),
    .Y(_03070_));
 sky130_fd_sc_hd__o21ba_1 _12279_ (.A1(_02899_),
    .A2(_02902_),
    .B1_N(_02900_),
    .X(_03071_));
 sky130_fd_sc_hd__and2b_2 _12280_ (.A_N(_03071_),
    .B(_03070_),
    .X(_03072_));
 sky130_fd_sc_hd__xnor2_1 _12281_ (.A(_03070_),
    .B(_03071_),
    .Y(_03073_));
 sky130_fd_sc_hd__and2_2 _12282_ (.A(_03065_),
    .B(_03073_),
    .X(_03074_));
 sky130_fd_sc_hd__nor2_1 _12283_ (.A(_03065_),
    .B(_03073_),
    .Y(_03075_));
 sky130_fd_sc_hd__or2_2 _12284_ (.A(_03074_),
    .B(_03075_),
    .X(_03076_));
 sky130_fd_sc_hd__a21o_4 _12285_ (.A1(_02885_),
    .A2(_02888_),
    .B1(_03076_),
    .X(_03077_));
 sky130_fd_sc_hd__nand3_2 _12286_ (.A(_02885_),
    .B(_02888_),
    .C(_03076_),
    .Y(_03078_));
 sky130_fd_sc_hd__o211ai_4 _12287_ (.A1(_02905_),
    .A2(_02907_),
    .B1(_03077_),
    .C1(_03078_),
    .Y(_03079_));
 sky130_fd_sc_hd__a211o_2 _12288_ (.A1(_03077_),
    .A2(_03078_),
    .B1(_02905_),
    .C1(_02907_),
    .X(_03080_));
 sky130_fd_sc_hd__a2bb2oi_4 _12289_ (.A1_N(_03059_),
    .A2_N(_03060_),
    .B1(_03079_),
    .B2(_03080_),
    .Y(_03081_));
 sky130_fd_sc_hd__and4bb_4 _12290_ (.A_N(_03059_),
    .B_N(_03060_),
    .C(_03079_),
    .D(_03080_),
    .X(_03082_));
 sky130_fd_sc_hd__a211o_2 _12291_ (.A1(_02892_),
    .A2(_02915_),
    .B1(_03081_),
    .C1(_03082_),
    .X(_03083_));
 sky130_fd_sc_hd__o211ai_4 _12292_ (.A1(_03081_),
    .A2(_03082_),
    .B1(_02892_),
    .C1(_02915_),
    .Y(_03084_));
 sky130_fd_sc_hd__o21ai_4 _12293_ (.A1(_02934_),
    .A2(_02935_),
    .B1(_02937_),
    .Y(_03085_));
 sky130_fd_sc_hd__a22oi_1 _12294_ (.A1(net327),
    .A2(net852),
    .B1(net862),
    .B2(net325),
    .Y(_03086_));
 sky130_fd_sc_hd__and4_1 _12295_ (.A(net325),
    .B(net327),
    .C(net852),
    .D(net862),
    .X(_03087_));
 sky130_fd_sc_hd__or2_1 _12296_ (.A(_03086_),
    .B(_03087_),
    .X(_03088_));
 sky130_fd_sc_hd__nand2_1 _12297_ (.A(\cla_inst.in2[29] ),
    .B(net841),
    .Y(_03089_));
 sky130_fd_sc_hd__nor2_2 _12298_ (.A(_03088_),
    .B(_03089_),
    .Y(_03090_));
 sky130_fd_sc_hd__and2_1 _12299_ (.A(_03088_),
    .B(_03089_),
    .X(_03091_));
 sky130_fd_sc_hd__nor2_2 _12300_ (.A(_03090_),
    .B(_03091_),
    .Y(_03092_));
 sky130_fd_sc_hd__a31o_2 _12301_ (.A1(net526),
    .A2(net633),
    .A3(_02896_),
    .B1(_02895_),
    .X(_03093_));
 sky130_fd_sc_hd__and3_1 _12302_ (.A(net536),
    .B(net617),
    .C(_02722_),
    .X(_03094_));
 sky130_fd_sc_hd__xnor2_2 _12303_ (.A(_03093_),
    .B(_03094_),
    .Y(_03095_));
 sky130_fd_sc_hd__a21oi_2 _12304_ (.A1(_02930_),
    .A2(_02933_),
    .B1(_03095_),
    .Y(_03096_));
 sky130_fd_sc_hd__and3_1 _12305_ (.A(_02930_),
    .B(_02933_),
    .C(_03095_),
    .X(_03097_));
 sky130_fd_sc_hd__nor2_2 _12306_ (.A(_03096_),
    .B(_03097_),
    .Y(_03098_));
 sky130_fd_sc_hd__xnor2_2 _12307_ (.A(_03092_),
    .B(_03098_),
    .Y(_03099_));
 sky130_fd_sc_hd__a21oi_4 _12308_ (.A1(_02910_),
    .A2(_02912_),
    .B1(_03099_),
    .Y(_03100_));
 sky130_fd_sc_hd__and3_1 _12309_ (.A(_02910_),
    .B(_02912_),
    .C(_03099_),
    .X(_03101_));
 sky130_fd_sc_hd__nor2_4 _12310_ (.A(_03100_),
    .B(_03101_),
    .Y(_03102_));
 sky130_fd_sc_hd__xor2_2 _12311_ (.A(_03085_),
    .B(_03102_),
    .X(_03103_));
 sky130_fd_sc_hd__nand3_2 _12312_ (.A(_03083_),
    .B(_03084_),
    .C(_03103_),
    .Y(_03104_));
 sky130_fd_sc_hd__a21o_1 _12313_ (.A1(_03083_),
    .A2(_03084_),
    .B1(_03103_),
    .X(_03105_));
 sky130_fd_sc_hd__nand2_2 _12314_ (.A(_03104_),
    .B(_03105_),
    .Y(_03106_));
 sky130_fd_sc_hd__a21o_4 _12315_ (.A1(_02916_),
    .A2(_02944_),
    .B1(_03106_),
    .X(_03107_));
 sky130_fd_sc_hd__nand3_2 _12316_ (.A(_02916_),
    .B(_02944_),
    .C(_03106_),
    .Y(_03108_));
 sky130_fd_sc_hd__o21ai_4 _12317_ (.A1(_02977_),
    .A2(_02978_),
    .B1(_02980_),
    .Y(_03109_));
 sky130_fd_sc_hd__o21ba_4 _12318_ (.A1(_02918_),
    .A2(_02941_),
    .B1_N(_02940_),
    .X(_03110_));
 sky130_fd_sc_hd__a22oi_4 _12319_ (.A1(net373),
    .A2(net789),
    .B1(net800),
    .B2(net364),
    .Y(_03111_));
 sky130_fd_sc_hd__and4_2 _12320_ (.A(net364),
    .B(net373),
    .C(net789),
    .D(net800),
    .X(_03112_));
 sky130_fd_sc_hd__nand2_1 _12321_ (.A(net383),
    .B(net778),
    .Y(_03113_));
 sky130_fd_sc_hd__o21a_1 _12322_ (.A1(_03111_),
    .A2(_03112_),
    .B1(_03113_),
    .X(_03114_));
 sky130_fd_sc_hd__nor3_2 _12323_ (.A(_03111_),
    .B(_03112_),
    .C(_03113_),
    .Y(_03115_));
 sky130_fd_sc_hd__nor2_1 _12324_ (.A(_03114_),
    .B(_03115_),
    .Y(_03116_));
 sky130_fd_sc_hd__or3_1 _12325_ (.A(_02951_),
    .B(_02954_),
    .C(_03116_),
    .X(_03117_));
 sky130_fd_sc_hd__o21ai_1 _12326_ (.A1(_02951_),
    .A2(_02954_),
    .B1(_03116_),
    .Y(_03118_));
 sky130_fd_sc_hd__and2_1 _12327_ (.A(_03117_),
    .B(_03118_),
    .X(_03119_));
 sky130_fd_sc_hd__nand3_2 _12328_ (.A(net389),
    .B(net766),
    .C(_03119_),
    .Y(_03120_));
 sky130_fd_sc_hd__a21o_1 _12329_ (.A1(net389),
    .A2(net766),
    .B1(_03119_),
    .X(_03121_));
 sky130_fd_sc_hd__nand2_2 _12330_ (.A(_03120_),
    .B(_03121_),
    .Y(_03122_));
 sky130_fd_sc_hd__inv_2 _12331_ (.A(_03122_),
    .Y(_03123_));
 sky130_fd_sc_hd__a31o_2 _12332_ (.A1(net388),
    .A2(net778),
    .A3(_02958_),
    .B1(_02957_),
    .X(_03124_));
 sky130_fd_sc_hd__xnor2_1 _12333_ (.A(_03122_),
    .B(_03124_),
    .Y(_03125_));
 sky130_fd_sc_hd__and3_2 _12334_ (.A(net396),
    .B(net755),
    .C(_03125_),
    .X(_03126_));
 sky130_fd_sc_hd__a21oi_2 _12335_ (.A1(net396),
    .A2(net755),
    .B1(_03125_),
    .Y(_03127_));
 sky130_fd_sc_hd__nor2_4 _12336_ (.A(_03126_),
    .B(_03127_),
    .Y(_03128_));
 sky130_fd_sc_hd__a22oi_2 _12337_ (.A1(net350),
    .A2(net821),
    .B1(net831),
    .B2(net342),
    .Y(_03129_));
 sky130_fd_sc_hd__and4_1 _12338_ (.A(net342),
    .B(net350),
    .C(net821),
    .D(net831),
    .X(_03130_));
 sky130_fd_sc_hd__nor2_1 _12339_ (.A(_03129_),
    .B(_03130_),
    .Y(_03131_));
 sky130_fd_sc_hd__nand2_2 _12340_ (.A(net358),
    .B(net810),
    .Y(_03132_));
 sky130_fd_sc_hd__xnor2_2 _12341_ (.A(_03131_),
    .B(_03132_),
    .Y(_03133_));
 sky130_fd_sc_hd__o21a_1 _12342_ (.A1(_02920_),
    .A2(_02923_),
    .B1(_03133_),
    .X(_03134_));
 sky130_fd_sc_hd__nor3_1 _12343_ (.A(_02920_),
    .B(_02923_),
    .C(_03133_),
    .Y(_03135_));
 sky130_fd_sc_hd__nor2_1 _12344_ (.A(_03134_),
    .B(_03135_),
    .Y(_03136_));
 sky130_fd_sc_hd__o21ba_1 _12345_ (.A1(_02966_),
    .A2(_02969_),
    .B1_N(_02967_),
    .X(_03137_));
 sky130_fd_sc_hd__xor2_1 _12346_ (.A(_03136_),
    .B(_03137_),
    .X(_03138_));
 sky130_fd_sc_hd__o21ba_1 _12347_ (.A1(_02972_),
    .A2(_02974_),
    .B1_N(_02971_),
    .X(_03139_));
 sky130_fd_sc_hd__or2_4 _12348_ (.A(_03138_),
    .B(_03139_),
    .X(_03140_));
 sky130_fd_sc_hd__nand2_1 _12349_ (.A(_03138_),
    .B(_03139_),
    .Y(_03141_));
 sky130_fd_sc_hd__and2_1 _12350_ (.A(_03140_),
    .B(_03141_),
    .X(_03142_));
 sky130_fd_sc_hd__or3b_1 _12351_ (.A(_02975_),
    .B(_02976_),
    .C_N(_03142_),
    .X(_03143_));
 sky130_fd_sc_hd__o21bai_1 _12352_ (.A1(_02975_),
    .A2(_02976_),
    .B1_N(_03142_),
    .Y(_03144_));
 sky130_fd_sc_hd__and2_2 _12353_ (.A(_03143_),
    .B(_03144_),
    .X(_03145_));
 sky130_fd_sc_hd__xnor2_4 _12354_ (.A(_03128_),
    .B(_03145_),
    .Y(_03146_));
 sky130_fd_sc_hd__xnor2_4 _12355_ (.A(_03110_),
    .B(_03146_),
    .Y(_03147_));
 sky130_fd_sc_hd__and2b_1 _12356_ (.A_N(_03147_),
    .B(_03109_),
    .X(_03148_));
 sky130_fd_sc_hd__xnor2_4 _12357_ (.A(_03109_),
    .B(_03147_),
    .Y(_03149_));
 sky130_fd_sc_hd__nand3_4 _12358_ (.A(_03107_),
    .B(_03108_),
    .C(_03149_),
    .Y(_03150_));
 sky130_fd_sc_hd__a21o_1 _12359_ (.A1(_03107_),
    .A2(_03108_),
    .B1(_03149_),
    .X(_03151_));
 sky130_fd_sc_hd__nand2_2 _12360_ (.A(_02946_),
    .B(_02986_),
    .Y(_03152_));
 sky130_fd_sc_hd__nand3_1 _12361_ (.A(_03150_),
    .B(_03151_),
    .C(_03152_),
    .Y(_03153_));
 sky130_fd_sc_hd__a21o_1 _12362_ (.A1(_03150_),
    .A2(_03151_),
    .B1(_03152_),
    .X(_03154_));
 sky130_fd_sc_hd__a31o_1 _12363_ (.A1(_02949_),
    .A2(_02980_),
    .A3(_02981_),
    .B1(_02984_),
    .X(_03155_));
 sky130_fd_sc_hd__and3_2 _12364_ (.A(_03153_),
    .B(_03154_),
    .C(_03155_),
    .X(_03156_));
 sky130_fd_sc_hd__a21oi_2 _12365_ (.A1(_03153_),
    .A2(_03154_),
    .B1(_03155_),
    .Y(_03157_));
 sky130_fd_sc_hd__or2_4 _12366_ (.A(_03156_),
    .B(_03157_),
    .X(_03158_));
 sky130_fd_sc_hd__and2b_4 _12367_ (.A_N(_02988_),
    .B(_02991_),
    .X(_03159_));
 sky130_fd_sc_hd__xnor2_4 _12368_ (.A(_03158_),
    .B(_03159_),
    .Y(_03160_));
 sky130_fd_sc_hd__o21ba_4 _12369_ (.A1(_02962_),
    .A2(_02964_),
    .B1_N(_02961_),
    .X(_03161_));
 sky130_fd_sc_hd__xnor2_4 _12370_ (.A(_03160_),
    .B(_03161_),
    .Y(_03162_));
 sky130_fd_sc_hd__nor2_4 _12371_ (.A(_02994_),
    .B(_02996_),
    .Y(_03163_));
 sky130_fd_sc_hd__or2_4 _12372_ (.A(_03162_),
    .B(_03163_),
    .X(_03164_));
 sky130_fd_sc_hd__xnor2_4 _12373_ (.A(_03162_),
    .B(_03163_),
    .Y(_03165_));
 sky130_fd_sc_hd__nand2_2 _12374_ (.A(_02808_),
    .B(_03001_),
    .Y(_03166_));
 sky130_fd_sc_hd__nor2_1 _12375_ (.A(_02806_),
    .B(_02999_),
    .Y(_03167_));
 sky130_fd_sc_hd__o22ai_4 _12376_ (.A1(_02809_),
    .A2(_03166_),
    .B1(_03167_),
    .B2(_03000_),
    .Y(_03168_));
 sky130_fd_sc_hd__nor2_2 _12377_ (.A(_02810_),
    .B(_03166_),
    .Y(_03169_));
 sky130_fd_sc_hd__a21oi_2 _12378_ (.A1(_02574_),
    .A2(_03169_),
    .B1(_03168_),
    .Y(_03170_));
 sky130_fd_sc_hd__or2_4 _12379_ (.A(_03165_),
    .B(_03170_),
    .X(_03171_));
 sky130_fd_sc_hd__nand2_1 _12380_ (.A(net260),
    .B(_03171_),
    .Y(_03172_));
 sky130_fd_sc_hd__a21o_2 _12381_ (.A1(_03165_),
    .A2(_03170_),
    .B1(_03172_),
    .X(_03173_));
 sky130_fd_sc_hd__mux2_1 _12382_ (.A0(_02836_),
    .A1(_02838_),
    .S(net291),
    .X(_03174_));
 sky130_fd_sc_hd__mux2_1 _12383_ (.A0(_02840_),
    .A1(_02843_),
    .S(net291),
    .X(_03175_));
 sky130_fd_sc_hd__mux2_1 _12384_ (.A0(_03174_),
    .A1(_03175_),
    .S(net296),
    .X(_03176_));
 sky130_fd_sc_hd__mux2_1 _12385_ (.A0(_02845_),
    .A1(_02847_),
    .S(net291),
    .X(_03177_));
 sky130_fd_sc_hd__mux2_1 _12386_ (.A0(_02814_),
    .A1(_02849_),
    .S(net597),
    .X(_03178_));
 sky130_fd_sc_hd__mux2_1 _12387_ (.A0(_03177_),
    .A1(_03178_),
    .S(net296),
    .X(_03179_));
 sky130_fd_sc_hd__mux2_1 _12388_ (.A0(_03176_),
    .A1(_03179_),
    .S(net301),
    .X(_03180_));
 sky130_fd_sc_hd__mux2_1 _12389_ (.A0(_02816_),
    .A1(_02818_),
    .S(net290),
    .X(_03181_));
 sky130_fd_sc_hd__mux2_1 _12390_ (.A0(_02820_),
    .A1(_02825_),
    .S(net287),
    .X(_03183_));
 sky130_fd_sc_hd__mux2_1 _12391_ (.A0(_03181_),
    .A1(_03183_),
    .S(net295),
    .X(_03184_));
 sky130_fd_sc_hd__mux2_2 _12392_ (.A0(_02823_),
    .A1(_02827_),
    .S(net596),
    .X(_03185_));
 sky130_fd_sc_hd__nor2_2 _12393_ (.A(net295),
    .B(_03185_),
    .Y(_03186_));
 sky130_fd_sc_hd__inv_2 _12394_ (.A(_03186_),
    .Y(_03187_));
 sky130_fd_sc_hd__mux2_1 _12395_ (.A0(_03184_),
    .A1(_03187_),
    .S(net301),
    .X(_03188_));
 sky130_fd_sc_hd__mux2_1 _12396_ (.A0(_03180_),
    .A1(_03188_),
    .S(net305),
    .X(_03189_));
 sky130_fd_sc_hd__or2_1 _12397_ (.A(net597),
    .B(_02853_),
    .X(_03190_));
 sky130_fd_sc_hd__mux2_1 _12398_ (.A0(_02834_),
    .A1(_02855_),
    .S(net597),
    .X(_03191_));
 sky130_fd_sc_hd__mux2_1 _12399_ (.A0(_03190_),
    .A1(_03191_),
    .S(net296),
    .X(_03192_));
 sky130_fd_sc_hd__or2_2 _12400_ (.A(net568),
    .B(_03192_),
    .X(_03194_));
 sky130_fd_sc_hd__or2_1 _12401_ (.A(net206),
    .B(_03194_),
    .X(_03195_));
 sky130_fd_sc_hd__a22o_1 _12402_ (.A1(_03193_),
    .A2(_03189_),
    .B1(_03195_),
    .B2(net208),
    .X(_03196_));
 sky130_fd_sc_hd__nand2_1 _12403_ (.A(_03173_),
    .B(_03196_),
    .Y(_08677_));
 sky130_fd_sc_hd__a22oi_1 _12404_ (.A1(net426),
    .A2(net725),
    .B1(net742),
    .B2(net410),
    .Y(_03197_));
 sky130_fd_sc_hd__and4_2 _12405_ (.A(net410),
    .B(net426),
    .C(net725),
    .D(net742),
    .X(_03198_));
 sky130_fd_sc_hd__nor2_1 _12406_ (.A(_03197_),
    .B(_03198_),
    .Y(_03199_));
 sky130_fd_sc_hd__a21oi_2 _12407_ (.A1(net417),
    .A2(net733),
    .B1(_03199_),
    .Y(_03200_));
 sky130_fd_sc_hd__and3_4 _12408_ (.A(net417),
    .B(net733),
    .C(_03199_),
    .X(_03201_));
 sky130_fd_sc_hd__nor2_4 _12409_ (.A(_03200_),
    .B(_03201_),
    .Y(_03202_));
 sky130_fd_sc_hd__a31o_4 _12410_ (.A1(net417),
    .A2(net742),
    .A3(_03028_),
    .B1(_03027_),
    .X(_03204_));
 sky130_fd_sc_hd__and2_1 _12411_ (.A(_03202_),
    .B(_03204_),
    .X(_03205_));
 sky130_fd_sc_hd__xor2_4 _12412_ (.A(_03202_),
    .B(_03204_),
    .X(_03206_));
 sky130_fd_sc_hd__a22oi_4 _12413_ (.A1(net444),
    .A2(net706),
    .B1(net715),
    .B2(net433),
    .Y(_03207_));
 sky130_fd_sc_hd__and4_1 _12414_ (.A(net433),
    .B(net444),
    .C(net706),
    .D(net715),
    .X(_03208_));
 sky130_fd_sc_hd__nor2_2 _12415_ (.A(_03207_),
    .B(_03208_),
    .Y(_03209_));
 sky130_fd_sc_hd__nand2_4 _12416_ (.A(net450),
    .B(net699),
    .Y(_03210_));
 sky130_fd_sc_hd__xnor2_4 _12417_ (.A(_03209_),
    .B(_03210_),
    .Y(_03211_));
 sky130_fd_sc_hd__and2_1 _12418_ (.A(_03206_),
    .B(_03211_),
    .X(_03212_));
 sky130_fd_sc_hd__xnor2_4 _12419_ (.A(_03206_),
    .B(_03211_),
    .Y(_03213_));
 sky130_fd_sc_hd__a21o_4 _12420_ (.A1(_03032_),
    .A2(_03041_),
    .B1(_03213_),
    .X(_03215_));
 sky130_fd_sc_hd__nand3_4 _12421_ (.A(_03032_),
    .B(_03041_),
    .C(_03213_),
    .Y(_03216_));
 sky130_fd_sc_hd__o21ba_4 _12422_ (.A1(_03047_),
    .A2(_03050_),
    .B1_N(_03048_),
    .X(_03217_));
 sky130_fd_sc_hd__a22oi_2 _12423_ (.A1(net465),
    .A2(net678),
    .B1(net686),
    .B2(net455),
    .Y(_03218_));
 sky130_fd_sc_hd__and4_1 _12424_ (.A(net455),
    .B(net465),
    .C(net678),
    .D(net686),
    .X(_03219_));
 sky130_fd_sc_hd__nor2_1 _12425_ (.A(_03218_),
    .B(_03219_),
    .Y(_03220_));
 sky130_fd_sc_hd__nand2_2 _12426_ (.A(net479),
    .B(net668),
    .Y(_03221_));
 sky130_fd_sc_hd__xnor2_2 _12427_ (.A(_03220_),
    .B(_03221_),
    .Y(_03222_));
 sky130_fd_sc_hd__o21a_4 _12428_ (.A1(_03035_),
    .A2(_03038_),
    .B1(_03222_),
    .X(_03223_));
 sky130_fd_sc_hd__nor3_2 _12429_ (.A(_03035_),
    .B(_03038_),
    .C(_03222_),
    .Y(_03224_));
 sky130_fd_sc_hd__nor2_4 _12430_ (.A(_03223_),
    .B(_03224_),
    .Y(_03226_));
 sky130_fd_sc_hd__and2b_1 _12431_ (.A_N(_03217_),
    .B(_03226_),
    .X(_03227_));
 sky130_fd_sc_hd__xnor2_4 _12432_ (.A(_03217_),
    .B(_03226_),
    .Y(_03228_));
 sky130_fd_sc_hd__a21o_1 _12433_ (.A1(_03215_),
    .A2(_03216_),
    .B1(_03228_),
    .X(_03229_));
 sky130_fd_sc_hd__nand3_4 _12434_ (.A(_03215_),
    .B(_03216_),
    .C(_03228_),
    .Y(_03230_));
 sky130_fd_sc_hd__nand2_2 _12435_ (.A(_03229_),
    .B(_03230_),
    .Y(_03231_));
 sky130_fd_sc_hd__a21o_4 _12436_ (.A1(_03043_),
    .A2(_03057_),
    .B1(_03231_),
    .X(_03232_));
 sky130_fd_sc_hd__nand3_4 _12437_ (.A(_03043_),
    .B(_03057_),
    .C(_03231_),
    .Y(_03233_));
 sky130_fd_sc_hd__a22oi_1 _12438_ (.A1(net519),
    .A2(net626),
    .B1(net634),
    .B2(net511),
    .Y(_03234_));
 sky130_fd_sc_hd__and4_1 _12439_ (.A(net511),
    .B(net519),
    .C(net626),
    .D(net634),
    .X(_03235_));
 sky130_fd_sc_hd__nor2_1 _12440_ (.A(_03234_),
    .B(_03235_),
    .Y(_03237_));
 sky130_fd_sc_hd__a21oi_2 _12441_ (.A1(net528),
    .A2(net617),
    .B1(_03237_),
    .Y(_03238_));
 sky130_fd_sc_hd__and3_2 _12442_ (.A(net528),
    .B(net618),
    .C(_03237_),
    .X(_03239_));
 sky130_fd_sc_hd__nor2_4 _12443_ (.A(_03238_),
    .B(_03239_),
    .Y(_03240_));
 sky130_fd_sc_hd__a22oi_4 _12444_ (.A1(net494),
    .A2(net655),
    .B1(net663),
    .B2(net484),
    .Y(_03241_));
 sky130_fd_sc_hd__and4_1 _12445_ (.A(net484),
    .B(net494),
    .C(net655),
    .D(net663),
    .X(_03242_));
 sky130_fd_sc_hd__nor2_2 _12446_ (.A(_03241_),
    .B(_03242_),
    .Y(_03243_));
 sky130_fd_sc_hd__nand2_4 _12447_ (.A(net503),
    .B(net645),
    .Y(_03244_));
 sky130_fd_sc_hd__xnor2_4 _12448_ (.A(_03243_),
    .B(_03244_),
    .Y(_03245_));
 sky130_fd_sc_hd__o21ba_2 _12449_ (.A1(_03066_),
    .A2(_03069_),
    .B1_N(_03067_),
    .X(_03246_));
 sky130_fd_sc_hd__and2b_1 _12450_ (.A_N(_03246_),
    .B(_03245_),
    .X(_03248_));
 sky130_fd_sc_hd__xnor2_4 _12451_ (.A(_03245_),
    .B(_03246_),
    .Y(_03249_));
 sky130_fd_sc_hd__xnor2_2 _12452_ (.A(_03240_),
    .B(_03249_),
    .Y(_03250_));
 sky130_fd_sc_hd__a21o_2 _12453_ (.A1(_03052_),
    .A2(_03054_),
    .B1(_03250_),
    .X(_03251_));
 sky130_fd_sc_hd__nand3_2 _12454_ (.A(_03052_),
    .B(_03054_),
    .C(_03250_),
    .Y(_03252_));
 sky130_fd_sc_hd__o211ai_4 _12455_ (.A1(_03072_),
    .A2(_03074_),
    .B1(_03251_),
    .C1(_03252_),
    .Y(_03253_));
 sky130_fd_sc_hd__a211o_2 _12456_ (.A1(_03251_),
    .A2(_03252_),
    .B1(_03072_),
    .C1(_03074_),
    .X(_03254_));
 sky130_fd_sc_hd__a22o_2 _12457_ (.A1(_03232_),
    .A2(_03233_),
    .B1(_03253_),
    .B2(_03254_),
    .X(_03255_));
 sky130_fd_sc_hd__nand4_4 _12458_ (.A(_03232_),
    .B(_03233_),
    .C(_03253_),
    .D(_03254_),
    .Y(_03256_));
 sky130_fd_sc_hd__o211ai_4 _12459_ (.A1(_03059_),
    .A2(_03082_),
    .B1(_03255_),
    .C1(_03256_),
    .Y(_03257_));
 sky130_fd_sc_hd__a211o_2 _12460_ (.A1(_03255_),
    .A2(_03256_),
    .B1(_03059_),
    .C1(_03082_),
    .X(_03259_));
 sky130_fd_sc_hd__a21o_4 _12461_ (.A1(_03092_),
    .A2(_03098_),
    .B1(_03096_),
    .X(_03260_));
 sky130_fd_sc_hd__a22oi_1 _12462_ (.A1(net327),
    .A2(net841),
    .B1(net852),
    .B2(net325),
    .Y(_03261_));
 sky130_fd_sc_hd__and4_1 _12463_ (.A(net325),
    .B(net327),
    .C(net841),
    .D(net852),
    .X(_03262_));
 sky130_fd_sc_hd__or2_1 _12464_ (.A(_03261_),
    .B(_03262_),
    .X(_03263_));
 sky130_fd_sc_hd__nand2_1 _12465_ (.A(net335),
    .B(net831),
    .Y(_03264_));
 sky130_fd_sc_hd__nor2_2 _12466_ (.A(_03263_),
    .B(_03264_),
    .Y(_03265_));
 sky130_fd_sc_hd__and2_1 _12467_ (.A(_03263_),
    .B(_03264_),
    .X(_03266_));
 sky130_fd_sc_hd__nor2_4 _12468_ (.A(_03265_),
    .B(_03266_),
    .Y(_03267_));
 sky130_fd_sc_hd__o21ba_4 _12469_ (.A1(_03061_),
    .A2(_03064_),
    .B1_N(_03062_),
    .X(_03268_));
 sky130_fd_sc_hd__nand2b_1 _12470_ (.A_N(_03093_),
    .B(_02722_),
    .Y(_03270_));
 sky130_fd_sc_hd__and3_4 _12471_ (.A(net549),
    .B(net617),
    .C(_03270_),
    .X(_03271_));
 sky130_fd_sc_hd__nand2b_1 _12472_ (.A_N(_03268_),
    .B(_03271_),
    .Y(_03272_));
 sky130_fd_sc_hd__xnor2_4 _12473_ (.A(_03268_),
    .B(_03271_),
    .Y(_03273_));
 sky130_fd_sc_hd__xnor2_4 _12474_ (.A(_03267_),
    .B(_03273_),
    .Y(_03274_));
 sky130_fd_sc_hd__a21oi_4 _12475_ (.A1(_03077_),
    .A2(_03079_),
    .B1(_03274_),
    .Y(_03275_));
 sky130_fd_sc_hd__and3_1 _12476_ (.A(_03077_),
    .B(_03079_),
    .C(_03274_),
    .X(_03276_));
 sky130_fd_sc_hd__nor2_4 _12477_ (.A(_03275_),
    .B(_03276_),
    .Y(_03277_));
 sky130_fd_sc_hd__xor2_4 _12478_ (.A(_03260_),
    .B(_03277_),
    .X(_03278_));
 sky130_fd_sc_hd__a21oi_2 _12479_ (.A1(_03257_),
    .A2(_03259_),
    .B1(_03278_),
    .Y(_03279_));
 sky130_fd_sc_hd__and3_1 _12480_ (.A(_03257_),
    .B(_03259_),
    .C(_03278_),
    .X(_03281_));
 sky130_fd_sc_hd__nand3_2 _12481_ (.A(_03257_),
    .B(_03259_),
    .C(_03278_),
    .Y(_03282_));
 sky130_fd_sc_hd__a211oi_2 _12482_ (.A1(_03083_),
    .A2(_03104_),
    .B1(_03279_),
    .C1(_03281_),
    .Y(_03283_));
 sky130_fd_sc_hd__o211a_1 _12483_ (.A1(_03279_),
    .A2(_03281_),
    .B1(_03083_),
    .C1(_03104_),
    .X(_03284_));
 sky130_fd_sc_hd__a21bo_2 _12484_ (.A1(_03128_),
    .A2(_03144_),
    .B1_N(_03143_),
    .X(_03285_));
 sky130_fd_sc_hd__a21oi_4 _12485_ (.A1(_03085_),
    .A2(_03102_),
    .B1(_03100_),
    .Y(_03286_));
 sky130_fd_sc_hd__a22oi_4 _12486_ (.A1(net373),
    .A2(net778),
    .B1(net789),
    .B2(net364),
    .Y(_03287_));
 sky130_fd_sc_hd__and4_4 _12487_ (.A(net364),
    .B(net373),
    .C(net778),
    .D(net789),
    .X(_03288_));
 sky130_fd_sc_hd__nand2_2 _12488_ (.A(net383),
    .B(net767),
    .Y(_03289_));
 sky130_fd_sc_hd__o21a_1 _12489_ (.A1(_03287_),
    .A2(_03288_),
    .B1(_03289_),
    .X(_03290_));
 sky130_fd_sc_hd__nor3_4 _12490_ (.A(_03287_),
    .B(_03288_),
    .C(_03289_),
    .Y(_03292_));
 sky130_fd_sc_hd__nor2_1 _12491_ (.A(_03290_),
    .B(_03292_),
    .Y(_03293_));
 sky130_fd_sc_hd__nor3_1 _12492_ (.A(_03112_),
    .B(_03115_),
    .C(_03293_),
    .Y(_03294_));
 sky130_fd_sc_hd__o21a_1 _12493_ (.A1(_03112_),
    .A2(_03115_),
    .B1(_03293_),
    .X(_03295_));
 sky130_fd_sc_hd__nor2_1 _12494_ (.A(_03294_),
    .B(_03295_),
    .Y(_03296_));
 sky130_fd_sc_hd__nand2_1 _12495_ (.A(net389),
    .B(net755),
    .Y(_03297_));
 sky130_fd_sc_hd__xor2_1 _12496_ (.A(_03296_),
    .B(_03297_),
    .X(_03298_));
 sky130_fd_sc_hd__a21oi_1 _12497_ (.A1(_03118_),
    .A2(_03120_),
    .B1(_03298_),
    .Y(_03299_));
 sky130_fd_sc_hd__and3_1 _12498_ (.A(_03118_),
    .B(_03120_),
    .C(_03298_),
    .X(_03300_));
 sky130_fd_sc_hd__nor2_2 _12499_ (.A(_03299_),
    .B(_03300_),
    .Y(_03301_));
 sky130_fd_sc_hd__nand2_4 _12500_ (.A(net399),
    .B(net746),
    .Y(_03303_));
 sky130_fd_sc_hd__xnor2_4 _12501_ (.A(_03301_),
    .B(_03303_),
    .Y(_03304_));
 sky130_fd_sc_hd__a22oi_2 _12502_ (.A1(net350),
    .A2(net812),
    .B1(net823),
    .B2(net342),
    .Y(_03305_));
 sky130_fd_sc_hd__and4_1 _12503_ (.A(net342),
    .B(net350),
    .C(net812),
    .D(net823),
    .X(_03306_));
 sky130_fd_sc_hd__nor2_1 _12504_ (.A(_03305_),
    .B(_03306_),
    .Y(_03307_));
 sky130_fd_sc_hd__nand2_2 _12505_ (.A(net358),
    .B(net800),
    .Y(_03308_));
 sky130_fd_sc_hd__xnor2_2 _12506_ (.A(_03307_),
    .B(_03308_),
    .Y(_03309_));
 sky130_fd_sc_hd__o21a_1 _12507_ (.A1(_03087_),
    .A2(_03090_),
    .B1(_03309_),
    .X(_03310_));
 sky130_fd_sc_hd__nor3_2 _12508_ (.A(_03087_),
    .B(_03090_),
    .C(_03309_),
    .Y(_03311_));
 sky130_fd_sc_hd__nor2_4 _12509_ (.A(_03310_),
    .B(_03311_),
    .Y(_03312_));
 sky130_fd_sc_hd__o21ba_2 _12510_ (.A1(_03129_),
    .A2(_03132_),
    .B1_N(_03130_),
    .X(_03314_));
 sky130_fd_sc_hd__xor2_4 _12511_ (.A(_03312_),
    .B(_03314_),
    .X(_03315_));
 sky130_fd_sc_hd__o21ba_2 _12512_ (.A1(_03135_),
    .A2(_03137_),
    .B1_N(_03134_),
    .X(_03316_));
 sky130_fd_sc_hd__nor2_4 _12513_ (.A(_03315_),
    .B(_03316_),
    .Y(_03317_));
 sky130_fd_sc_hd__and2_1 _12514_ (.A(_03315_),
    .B(_03316_),
    .X(_03318_));
 sky130_fd_sc_hd__nor2_4 _12515_ (.A(_03317_),
    .B(_03318_),
    .Y(_03319_));
 sky130_fd_sc_hd__nand2b_1 _12516_ (.A_N(_03140_),
    .B(_03319_),
    .Y(_03320_));
 sky130_fd_sc_hd__xnor2_4 _12517_ (.A(_03140_),
    .B(_03319_),
    .Y(_03321_));
 sky130_fd_sc_hd__xnor2_4 _12518_ (.A(_03304_),
    .B(_03321_),
    .Y(_03322_));
 sky130_fd_sc_hd__xnor2_2 _12519_ (.A(_03286_),
    .B(_03322_),
    .Y(_03323_));
 sky130_fd_sc_hd__nand2b_1 _12520_ (.A_N(_03323_),
    .B(_03285_),
    .Y(_03325_));
 sky130_fd_sc_hd__xor2_2 _12521_ (.A(_03285_),
    .B(_03323_),
    .X(_03326_));
 sky130_fd_sc_hd__or3_1 _12522_ (.A(_03283_),
    .B(_03284_),
    .C(_03326_),
    .X(_03327_));
 sky130_fd_sc_hd__o21ai_1 _12523_ (.A1(_03283_),
    .A2(_03284_),
    .B1(_03326_),
    .Y(_03328_));
 sky130_fd_sc_hd__nand2_2 _12524_ (.A(_03327_),
    .B(_03328_),
    .Y(_03329_));
 sky130_fd_sc_hd__a21oi_4 _12525_ (.A1(_03107_),
    .A2(_03150_),
    .B1(_03329_),
    .Y(_03330_));
 sky130_fd_sc_hd__and3_2 _12526_ (.A(_03107_),
    .B(_03150_),
    .C(_03329_),
    .X(_03331_));
 sky130_fd_sc_hd__o21ba_2 _12527_ (.A1(_03110_),
    .A2(_03146_),
    .B1_N(_03148_),
    .X(_03332_));
 sky130_fd_sc_hd__nor3_4 _12528_ (.A(_03330_),
    .B(_03331_),
    .C(_03332_),
    .Y(_03333_));
 sky130_fd_sc_hd__o21a_1 _12529_ (.A1(_03330_),
    .A2(_03331_),
    .B1(_03332_),
    .X(_03334_));
 sky130_fd_sc_hd__or2_4 _12530_ (.A(_03333_),
    .B(_03334_),
    .X(_03336_));
 sky130_fd_sc_hd__a31o_4 _12531_ (.A1(_03150_),
    .A2(_03151_),
    .A3(_03152_),
    .B1(_03156_),
    .X(_03337_));
 sky130_fd_sc_hd__nand2b_1 _12532_ (.A_N(_03336_),
    .B(_03337_),
    .Y(_03338_));
 sky130_fd_sc_hd__and2b_1 _12533_ (.A_N(_03337_),
    .B(_03336_),
    .X(_03339_));
 sky130_fd_sc_hd__xnor2_4 _12534_ (.A(_03336_),
    .B(_03337_),
    .Y(_03340_));
 sky130_fd_sc_hd__a21oi_4 _12535_ (.A1(_03123_),
    .A2(_03124_),
    .B1(_03126_),
    .Y(_03341_));
 sky130_fd_sc_hd__xnor2_4 _12536_ (.A(_03340_),
    .B(_03341_),
    .Y(_03342_));
 sky130_fd_sc_hd__o32ai_4 _12537_ (.A1(_03156_),
    .A2(_03157_),
    .A3(_03159_),
    .B1(_03160_),
    .B2(_03161_),
    .Y(_03343_));
 sky130_fd_sc_hd__nand2_1 _12538_ (.A(_03342_),
    .B(net116),
    .Y(_03344_));
 sky130_fd_sc_hd__nor2_1 _12539_ (.A(_03342_),
    .B(net116),
    .Y(_03345_));
 sky130_fd_sc_hd__xnor2_4 _12540_ (.A(_03342_),
    .B(net116),
    .Y(_03347_));
 sky130_fd_sc_hd__a21oi_2 _12541_ (.A1(_03164_),
    .A2(_03171_),
    .B1(_03347_),
    .Y(_03348_));
 sky130_fd_sc_hd__a311oi_4 _12542_ (.A1(_03164_),
    .A2(_03171_),
    .A3(_03347_),
    .B1(_03348_),
    .C1(net255),
    .Y(_03349_));
 sky130_fd_sc_hd__mux2_1 _12543_ (.A0(_02627_),
    .A1(_02633_),
    .S(net293),
    .X(_03350_));
 sky130_fd_sc_hd__mux2_1 _12544_ (.A0(_02600_),
    .A1(_02638_),
    .S(net586),
    .X(_03351_));
 sky130_fd_sc_hd__mux2_1 _12545_ (.A0(_03350_),
    .A1(_03351_),
    .S(net302),
    .X(_03352_));
 sky130_fd_sc_hd__and3_2 _12546_ (.A(net583),
    .B(net598),
    .C(_02607_),
    .X(_03353_));
 sky130_fd_sc_hd__mux2_1 _12547_ (.A0(_02605_),
    .A1(_02612_),
    .S(net293),
    .X(_03354_));
 sky130_fd_sc_hd__nor2_1 _12548_ (.A(net567),
    .B(_03353_),
    .Y(_03355_));
 sky130_fd_sc_hd__a21o_1 _12549_ (.A1(net567),
    .A2(_03354_),
    .B1(_03355_),
    .X(_03356_));
 sky130_fd_sc_hd__mux2_1 _12550_ (.A0(_03352_),
    .A1(_03356_),
    .S(net307),
    .X(_03358_));
 sky130_fd_sc_hd__mux2_1 _12551_ (.A0(_02622_),
    .A1(_02647_),
    .S(net586),
    .X(_03359_));
 sky130_fd_sc_hd__or2_2 _12552_ (.A(net567),
    .B(_03359_),
    .X(_03360_));
 sky130_fd_sc_hd__or2_1 _12553_ (.A(net206),
    .B(_03360_),
    .X(_03361_));
 sky130_fd_sc_hd__a22o_1 _12554_ (.A1(_03193_),
    .A2(_03358_),
    .B1(_03361_),
    .B2(net209),
    .X(_03362_));
 sky130_fd_sc_hd__nand2b_1 _12555_ (.A_N(_03349_),
    .B(_03362_),
    .Y(_08678_));
 sky130_fd_sc_hd__nand2_8 _12556_ (.A(net417),
    .B(net727),
    .Y(_03363_));
 sky130_fd_sc_hd__a22o_1 _12557_ (.A1(net423),
    .A2(net715),
    .B1(net733),
    .B2(net410),
    .X(_03364_));
 sky130_fd_sc_hd__and2_4 _12558_ (.A(net407),
    .B(net715),
    .X(_03365_));
 sky130_fd_sc_hd__a21bo_2 _12559_ (.A1(_03025_),
    .A2(_03365_),
    .B1_N(_03364_),
    .X(_03366_));
 sky130_fd_sc_hd__xor2_4 _12560_ (.A(_03363_),
    .B(_03366_),
    .X(_03368_));
 sky130_fd_sc_hd__or3_1 _12561_ (.A(_03198_),
    .B(_03201_),
    .C(_03368_),
    .X(_03369_));
 sky130_fd_sc_hd__o21ai_4 _12562_ (.A1(_03198_),
    .A2(_03201_),
    .B1(_03368_),
    .Y(_03370_));
 sky130_fd_sc_hd__and2_2 _12563_ (.A(_03369_),
    .B(_03370_),
    .X(_03371_));
 sky130_fd_sc_hd__a22oi_4 _12564_ (.A1(net442),
    .A2(net699),
    .B1(net706),
    .B2(net433),
    .Y(_03372_));
 sky130_fd_sc_hd__and4_1 _12565_ (.A(net433),
    .B(net442),
    .C(net699),
    .D(net706),
    .X(_03373_));
 sky130_fd_sc_hd__nor2_2 _12566_ (.A(_03372_),
    .B(_03373_),
    .Y(_03374_));
 sky130_fd_sc_hd__nand2_4 _12567_ (.A(net453),
    .B(net689),
    .Y(_03375_));
 sky130_fd_sc_hd__xnor2_4 _12568_ (.A(_03374_),
    .B(_03375_),
    .Y(_03376_));
 sky130_fd_sc_hd__nand2_1 _12569_ (.A(_03371_),
    .B(_03376_),
    .Y(_03377_));
 sky130_fd_sc_hd__xor2_2 _12570_ (.A(_03371_),
    .B(_03376_),
    .X(_03378_));
 sky130_fd_sc_hd__o21ai_2 _12571_ (.A1(_03205_),
    .A2(_03212_),
    .B1(_03378_),
    .Y(_03379_));
 sky130_fd_sc_hd__or3_2 _12572_ (.A(_03205_),
    .B(_03212_),
    .C(_03378_),
    .X(_03380_));
 sky130_fd_sc_hd__o21ba_2 _12573_ (.A1(_03218_),
    .A2(_03221_),
    .B1_N(_03219_),
    .X(_03381_));
 sky130_fd_sc_hd__o21ba_1 _12574_ (.A1(_03207_),
    .A2(_03210_),
    .B1_N(_03208_),
    .X(_03382_));
 sky130_fd_sc_hd__a22oi_4 _12575_ (.A1(net469),
    .A2(net671),
    .B1(net684),
    .B2(net460),
    .Y(_03383_));
 sky130_fd_sc_hd__and4_1 _12576_ (.A(net460),
    .B(net469),
    .C(net671),
    .D(net684),
    .X(_03384_));
 sky130_fd_sc_hd__nor2_1 _12577_ (.A(_03383_),
    .B(_03384_),
    .Y(_03385_));
 sky130_fd_sc_hd__nand2_2 _12578_ (.A(net479),
    .B(net663),
    .Y(_03386_));
 sky130_fd_sc_hd__xnor2_2 _12579_ (.A(_03385_),
    .B(_03386_),
    .Y(_03387_));
 sky130_fd_sc_hd__and2b_1 _12580_ (.A_N(_03382_),
    .B(_03387_),
    .X(_03389_));
 sky130_fd_sc_hd__xnor2_2 _12581_ (.A(_03382_),
    .B(_03387_),
    .Y(_03390_));
 sky130_fd_sc_hd__and2b_1 _12582_ (.A_N(_03381_),
    .B(_03390_),
    .X(_03391_));
 sky130_fd_sc_hd__xnor2_2 _12583_ (.A(_03381_),
    .B(_03390_),
    .Y(_03392_));
 sky130_fd_sc_hd__a21oi_1 _12584_ (.A1(_03379_),
    .A2(_03380_),
    .B1(_03392_),
    .Y(_03393_));
 sky130_fd_sc_hd__and3_1 _12585_ (.A(_03379_),
    .B(_03380_),
    .C(_03392_),
    .X(_03394_));
 sky130_fd_sc_hd__or2_4 _12586_ (.A(_03393_),
    .B(_03394_),
    .X(_03395_));
 sky130_fd_sc_hd__a21oi_4 _12587_ (.A1(_03215_),
    .A2(_03230_),
    .B1(_03395_),
    .Y(_03396_));
 sky130_fd_sc_hd__and3_2 _12588_ (.A(_03215_),
    .B(_03230_),
    .C(_03395_),
    .X(_03397_));
 sky130_fd_sc_hd__a21oi_4 _12589_ (.A1(_03240_),
    .A2(_03249_),
    .B1(_03248_),
    .Y(_03398_));
 sky130_fd_sc_hd__a22oi_1 _12590_ (.A1(net519),
    .A2(net617),
    .B1(net625),
    .B2(net511),
    .Y(_03400_));
 sky130_fd_sc_hd__nand2_1 _12591_ (.A(net511),
    .B(net619),
    .Y(_03401_));
 sky130_fd_sc_hd__and4_1 _12592_ (.A(net511),
    .B(net519),
    .C(net618),
    .D(net626),
    .X(_03402_));
 sky130_fd_sc_hd__or2_2 _12593_ (.A(_03400_),
    .B(_03402_),
    .X(_03403_));
 sky130_fd_sc_hd__a22oi_1 _12594_ (.A1(net495),
    .A2(net645),
    .B1(net655),
    .B2(net485),
    .Y(_03404_));
 sky130_fd_sc_hd__and4_2 _12595_ (.A(net484),
    .B(net494),
    .C(net645),
    .D(net655),
    .X(_03405_));
 sky130_fd_sc_hd__nor2_1 _12596_ (.A(_03404_),
    .B(_03405_),
    .Y(_03406_));
 sky130_fd_sc_hd__and2_1 _12597_ (.A(net503),
    .B(net635),
    .X(_03407_));
 sky130_fd_sc_hd__nor2_1 _12598_ (.A(_03406_),
    .B(_03407_),
    .Y(_03408_));
 sky130_fd_sc_hd__and2_2 _12599_ (.A(_03406_),
    .B(_03407_),
    .X(_03409_));
 sky130_fd_sc_hd__nor2_4 _12600_ (.A(_03408_),
    .B(_03409_),
    .Y(_03410_));
 sky130_fd_sc_hd__o21ba_2 _12601_ (.A1(_03241_),
    .A2(_03244_),
    .B1_N(_03242_),
    .X(_03411_));
 sky130_fd_sc_hd__nand2b_2 _12602_ (.A_N(_03411_),
    .B(_03410_),
    .Y(_03412_));
 sky130_fd_sc_hd__xnor2_4 _12603_ (.A(_03410_),
    .B(_03411_),
    .Y(_03413_));
 sky130_fd_sc_hd__nand2b_2 _12604_ (.A_N(_03403_),
    .B(_03413_),
    .Y(_03414_));
 sky130_fd_sc_hd__xnor2_2 _12605_ (.A(_03403_),
    .B(_03413_),
    .Y(_03415_));
 sky130_fd_sc_hd__o21ai_2 _12606_ (.A1(_03223_),
    .A2(_03227_),
    .B1(_03415_),
    .Y(_03416_));
 sky130_fd_sc_hd__or3_1 _12607_ (.A(_03223_),
    .B(_03227_),
    .C(_03415_),
    .X(_03417_));
 sky130_fd_sc_hd__nand2_2 _12608_ (.A(_03416_),
    .B(_03417_),
    .Y(_03418_));
 sky130_fd_sc_hd__or2_1 _12609_ (.A(_03398_),
    .B(_03418_),
    .X(_03419_));
 sky130_fd_sc_hd__xnor2_4 _12610_ (.A(_03398_),
    .B(_03418_),
    .Y(_03421_));
 sky130_fd_sc_hd__o21a_2 _12611_ (.A1(_03396_),
    .A2(_03397_),
    .B1(_03421_),
    .X(_03422_));
 sky130_fd_sc_hd__nor3_4 _12612_ (.A(_03396_),
    .B(_03397_),
    .C(_03421_),
    .Y(_03423_));
 sky130_fd_sc_hd__a211oi_4 _12613_ (.A1(_03232_),
    .A2(_03256_),
    .B1(_03422_),
    .C1(_03423_),
    .Y(_03424_));
 sky130_fd_sc_hd__o211a_2 _12614_ (.A1(_03422_),
    .A2(_03423_),
    .B1(_03232_),
    .C1(_03256_),
    .X(_03425_));
 sky130_fd_sc_hd__a21bo_4 _12615_ (.A1(_03267_),
    .A2(_03273_),
    .B1_N(_03272_),
    .X(_03426_));
 sky130_fd_sc_hd__or2_2 _12616_ (.A(_03235_),
    .B(_03239_),
    .X(_03427_));
 sky130_fd_sc_hd__a22oi_4 _12617_ (.A1(net328),
    .A2(net831),
    .B1(net841),
    .B2(net318),
    .Y(_03428_));
 sky130_fd_sc_hd__and4_1 _12618_ (.A(net318),
    .B(net328),
    .C(net831),
    .D(net841),
    .X(_03429_));
 sky130_fd_sc_hd__nor2_1 _12619_ (.A(_03428_),
    .B(_03429_),
    .Y(_03430_));
 sky130_fd_sc_hd__nand2_2 _12620_ (.A(net337),
    .B(net823),
    .Y(_03432_));
 sky130_fd_sc_hd__xnor2_2 _12621_ (.A(_03430_),
    .B(_03432_),
    .Y(_03433_));
 sky130_fd_sc_hd__nand2_4 _12622_ (.A(_03427_),
    .B(_03433_),
    .Y(_03434_));
 sky130_fd_sc_hd__or2_1 _12623_ (.A(_03427_),
    .B(_03433_),
    .X(_03435_));
 sky130_fd_sc_hd__nand2_1 _12624_ (.A(_03434_),
    .B(_03435_),
    .Y(_03436_));
 sky130_fd_sc_hd__a21o_2 _12625_ (.A1(_03251_),
    .A2(_03253_),
    .B1(_03436_),
    .X(_03437_));
 sky130_fd_sc_hd__nand3_1 _12626_ (.A(_03251_),
    .B(_03253_),
    .C(_03436_),
    .Y(_03438_));
 sky130_fd_sc_hd__nand2_2 _12627_ (.A(_03437_),
    .B(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__nand2b_1 _12628_ (.A_N(_03439_),
    .B(_03426_),
    .Y(_03440_));
 sky130_fd_sc_hd__xor2_4 _12629_ (.A(_03426_),
    .B(_03439_),
    .X(_03441_));
 sky130_fd_sc_hd__o21a_2 _12630_ (.A1(_03424_),
    .A2(_03425_),
    .B1(_03441_),
    .X(_03442_));
 sky130_fd_sc_hd__nor3_4 _12631_ (.A(_03424_),
    .B(_03425_),
    .C(_03441_),
    .Y(_03443_));
 sky130_fd_sc_hd__a211oi_4 _12632_ (.A1(_03257_),
    .A2(_03282_),
    .B1(_03442_),
    .C1(_03443_),
    .Y(_03444_));
 sky130_fd_sc_hd__o211a_1 _12633_ (.A1(_03442_),
    .A2(_03443_),
    .B1(_03257_),
    .C1(_03282_),
    .X(_03445_));
 sky130_fd_sc_hd__a21bo_2 _12634_ (.A1(_03304_),
    .A2(_03321_),
    .B1_N(_03320_),
    .X(_03446_));
 sky130_fd_sc_hd__a21oi_2 _12635_ (.A1(_03260_),
    .A2(_03277_),
    .B1(_03275_),
    .Y(_03447_));
 sky130_fd_sc_hd__a22oi_4 _12636_ (.A1(net376),
    .A2(net767),
    .B1(net778),
    .B2(net367),
    .Y(_03448_));
 sky130_fd_sc_hd__and4_2 _12637_ (.A(net367),
    .B(net376),
    .C(net767),
    .D(net778),
    .X(_03449_));
 sky130_fd_sc_hd__nand2_1 _12638_ (.A(net384),
    .B(net756),
    .Y(_03450_));
 sky130_fd_sc_hd__o21a_1 _12639_ (.A1(_03448_),
    .A2(_03449_),
    .B1(_03450_),
    .X(_03451_));
 sky130_fd_sc_hd__nor3_2 _12640_ (.A(_03448_),
    .B(_03449_),
    .C(_03450_),
    .Y(_03453_));
 sky130_fd_sc_hd__nor2_2 _12641_ (.A(_03451_),
    .B(_03453_),
    .Y(_03454_));
 sky130_fd_sc_hd__or3_1 _12642_ (.A(_03288_),
    .B(_03292_),
    .C(_03454_),
    .X(_03455_));
 sky130_fd_sc_hd__o21ai_4 _12643_ (.A1(_03288_),
    .A2(_03292_),
    .B1(_03454_),
    .Y(_03456_));
 sky130_fd_sc_hd__and2_2 _12644_ (.A(_03455_),
    .B(_03456_),
    .X(_03457_));
 sky130_fd_sc_hd__nand3_4 _12645_ (.A(net389),
    .B(net747),
    .C(_03457_),
    .Y(_03458_));
 sky130_fd_sc_hd__a21o_1 _12646_ (.A1(net389),
    .A2(net747),
    .B1(_03457_),
    .X(_03459_));
 sky130_fd_sc_hd__nand2_1 _12647_ (.A(_03458_),
    .B(_03459_),
    .Y(_03460_));
 sky130_fd_sc_hd__a31o_2 _12648_ (.A1(net389),
    .A2(net755),
    .A3(_03296_),
    .B1(_03295_),
    .X(_03461_));
 sky130_fd_sc_hd__nand2b_4 _12649_ (.A_N(_03460_),
    .B(_03461_),
    .Y(_03462_));
 sky130_fd_sc_hd__nand2b_1 _12650_ (.A_N(_03461_),
    .B(_03460_),
    .Y(_03464_));
 sky130_fd_sc_hd__nand2_1 _12651_ (.A(_03462_),
    .B(_03464_),
    .Y(_03465_));
 sky130_fd_sc_hd__nand2_1 _12652_ (.A(net399),
    .B(net738),
    .Y(_03466_));
 sky130_fd_sc_hd__or2_4 _12653_ (.A(_03465_),
    .B(_03466_),
    .X(_03467_));
 sky130_fd_sc_hd__nand2_1 _12654_ (.A(_03465_),
    .B(_03466_),
    .Y(_03468_));
 sky130_fd_sc_hd__and2_1 _12655_ (.A(_03467_),
    .B(_03468_),
    .X(_03469_));
 sky130_fd_sc_hd__a22oi_2 _12656_ (.A1(net350),
    .A2(net802),
    .B1(net812),
    .B2(net342),
    .Y(_03470_));
 sky130_fd_sc_hd__and4_1 _12657_ (.A(net342),
    .B(net350),
    .C(net802),
    .D(net812),
    .X(_03471_));
 sky130_fd_sc_hd__nor2_1 _12658_ (.A(_03470_),
    .B(_03471_),
    .Y(_03472_));
 sky130_fd_sc_hd__nand2_2 _12659_ (.A(net357),
    .B(net795),
    .Y(_03473_));
 sky130_fd_sc_hd__xnor2_2 _12660_ (.A(_03472_),
    .B(_03473_),
    .Y(_03474_));
 sky130_fd_sc_hd__o21a_1 _12661_ (.A1(_03262_),
    .A2(_03265_),
    .B1(_03474_),
    .X(_03475_));
 sky130_fd_sc_hd__nor3_2 _12662_ (.A(_03262_),
    .B(_03265_),
    .C(_03474_),
    .Y(_03476_));
 sky130_fd_sc_hd__nor2_1 _12663_ (.A(_03475_),
    .B(_03476_),
    .Y(_03477_));
 sky130_fd_sc_hd__o21ba_2 _12664_ (.A1(_03305_),
    .A2(_03308_),
    .B1_N(_03306_),
    .X(_03478_));
 sky130_fd_sc_hd__xor2_1 _12665_ (.A(_03477_),
    .B(_03478_),
    .X(_03479_));
 sky130_fd_sc_hd__o21ba_1 _12666_ (.A1(_03311_),
    .A2(_03314_),
    .B1_N(_03310_),
    .X(_03480_));
 sky130_fd_sc_hd__or2_2 _12667_ (.A(_03479_),
    .B(_03480_),
    .X(_03481_));
 sky130_fd_sc_hd__nand2_1 _12668_ (.A(_03479_),
    .B(_03480_),
    .Y(_03482_));
 sky130_fd_sc_hd__and2_2 _12669_ (.A(_03481_),
    .B(_03482_),
    .X(_03483_));
 sky130_fd_sc_hd__xor2_2 _12670_ (.A(_03317_),
    .B(_03483_),
    .X(_03485_));
 sky130_fd_sc_hd__xnor2_1 _12671_ (.A(_03469_),
    .B(_03485_),
    .Y(_03486_));
 sky130_fd_sc_hd__or2_2 _12672_ (.A(_03447_),
    .B(_03486_),
    .X(_03487_));
 sky130_fd_sc_hd__xnor2_1 _12673_ (.A(_03447_),
    .B(_03486_),
    .Y(_03488_));
 sky130_fd_sc_hd__nand2b_2 _12674_ (.A_N(_03488_),
    .B(_03446_),
    .Y(_03489_));
 sky130_fd_sc_hd__xor2_1 _12675_ (.A(_03446_),
    .B(_03488_),
    .X(_03490_));
 sky130_fd_sc_hd__or3_2 _12676_ (.A(_03444_),
    .B(_03445_),
    .C(_03490_),
    .X(_03491_));
 sky130_fd_sc_hd__inv_2 _12677_ (.A(_03491_),
    .Y(_03492_));
 sky130_fd_sc_hd__o21ai_1 _12678_ (.A1(_03444_),
    .A2(_03445_),
    .B1(_03490_),
    .Y(_03493_));
 sky130_fd_sc_hd__nand2_2 _12679_ (.A(_03491_),
    .B(_03493_),
    .Y(_03494_));
 sky130_fd_sc_hd__o21ba_1 _12680_ (.A1(_03284_),
    .A2(_03326_),
    .B1_N(_03283_),
    .X(_03496_));
 sky130_fd_sc_hd__nor2_1 _12681_ (.A(_03494_),
    .B(_03496_),
    .Y(_03497_));
 sky130_fd_sc_hd__xnor2_2 _12682_ (.A(_03494_),
    .B(_03496_),
    .Y(_03498_));
 sky130_fd_sc_hd__o21a_1 _12683_ (.A1(_03286_),
    .A2(_03322_),
    .B1(_03325_),
    .X(_03499_));
 sky130_fd_sc_hd__or2_2 _12684_ (.A(_03498_),
    .B(_03499_),
    .X(_03500_));
 sky130_fd_sc_hd__nand2_2 _12685_ (.A(_03498_),
    .B(_03499_),
    .Y(_03501_));
 sky130_fd_sc_hd__o211a_4 _12686_ (.A1(_03330_),
    .A2(_03333_),
    .B1(_03500_),
    .C1(_03501_),
    .X(_03502_));
 sky130_fd_sc_hd__a211oi_4 _12687_ (.A1(_03500_),
    .A2(_03501_),
    .B1(_03330_),
    .C1(_03333_),
    .Y(_03503_));
 sky130_fd_sc_hd__o21ba_2 _12688_ (.A1(_03300_),
    .A2(_03303_),
    .B1_N(_03299_),
    .X(_03504_));
 sky130_fd_sc_hd__nor3_4 _12689_ (.A(_03502_),
    .B(_03503_),
    .C(_03504_),
    .Y(_03505_));
 sky130_fd_sc_hd__o21a_1 _12690_ (.A1(_03502_),
    .A2(_03503_),
    .B1(_03504_),
    .X(_03507_));
 sky130_fd_sc_hd__or2_4 _12691_ (.A(_03505_),
    .B(_03507_),
    .X(_03508_));
 sky130_fd_sc_hd__o21a_2 _12692_ (.A1(_03339_),
    .A2(_03341_),
    .B1(_03338_),
    .X(_03509_));
 sky130_fd_sc_hd__or2_2 _12693_ (.A(_03508_),
    .B(_03509_),
    .X(_03510_));
 sky130_fd_sc_hd__xnor2_4 _12694_ (.A(_03508_),
    .B(_03509_),
    .Y(_03511_));
 sky130_fd_sc_hd__a21o_1 _12695_ (.A1(_03164_),
    .A2(_03344_),
    .B1(_03345_),
    .X(_03512_));
 sky130_fd_sc_hd__or2_1 _12696_ (.A(_03165_),
    .B(_03347_),
    .X(_03513_));
 sky130_fd_sc_hd__o21a_2 _12697_ (.A1(_03170_),
    .A2(_03513_),
    .B1(_03512_),
    .X(_03514_));
 sky130_fd_sc_hd__nor2_1 _12698_ (.A(_03511_),
    .B(_03514_),
    .Y(_03515_));
 sky130_fd_sc_hd__a21o_1 _12699_ (.A1(_03511_),
    .A2(_03514_),
    .B1(net255),
    .X(_03516_));
 sky130_fd_sc_hd__and4_2 _12700_ (.A(net584),
    .B(net596),
    .C(_05899_),
    .D(net213),
    .X(_03518_));
 sky130_fd_sc_hd__inv_2 _12701_ (.A(_03518_),
    .Y(_03519_));
 sky130_fd_sc_hd__mux2_1 _12702_ (.A0(_02821_),
    .A1(_02828_),
    .S(net294),
    .X(_03520_));
 sky130_fd_sc_hd__mux2_1 _12703_ (.A0(_03519_),
    .A1(_03520_),
    .S(net566),
    .X(_03521_));
 sky130_fd_sc_hd__mux4_1 _12704_ (.A0(_02814_),
    .A1(_02816_),
    .A2(_02847_),
    .A3(_02849_),
    .S0(net290),
    .S1(net584),
    .X(_03522_));
 sky130_fd_sc_hd__mux4_2 _12705_ (.A0(_02838_),
    .A1(_02840_),
    .A2(_02843_),
    .A3(_02845_),
    .S0(net291),
    .S1(net296),
    .X(_03523_));
 sky130_fd_sc_hd__mux2_1 _12706_ (.A0(_03522_),
    .A1(_03523_),
    .S(net566),
    .X(_03524_));
 sky130_fd_sc_hd__mux2_1 _12707_ (.A0(_03521_),
    .A1(_03524_),
    .S(net554),
    .X(_03525_));
 sky130_fd_sc_hd__mux4_2 _12708_ (.A0(_02834_),
    .A1(_02836_),
    .A2(_02853_),
    .A3(_02855_),
    .S0(net291),
    .S1(net585),
    .X(_03526_));
 sky130_fd_sc_hd__or2_4 _12709_ (.A(net575),
    .B(_03526_),
    .X(_03527_));
 sky130_fd_sc_hd__or2_1 _12710_ (.A(net206),
    .B(_03527_),
    .X(_03529_));
 sky130_fd_sc_hd__a22o_1 _12711_ (.A1(_03193_),
    .A2(_03525_),
    .B1(_03529_),
    .B2(net209),
    .X(_03530_));
 sky130_fd_sc_hd__o21ai_1 _12712_ (.A1(_03515_),
    .A2(_03516_),
    .B1(_03530_),
    .Y(_08679_));
 sky130_fd_sc_hd__a22oi_2 _12713_ (.A1(net423),
    .A2(net706),
    .B1(net725),
    .B2(net407),
    .Y(_03531_));
 sky130_fd_sc_hd__and4_1 _12714_ (.A(net407),
    .B(net423),
    .C(net706),
    .D(net725),
    .X(_03532_));
 sky130_fd_sc_hd__nor2_1 _12715_ (.A(_03531_),
    .B(_03532_),
    .Y(_03533_));
 sky130_fd_sc_hd__nand2_1 _12716_ (.A(net416),
    .B(net715),
    .Y(_03534_));
 sky130_fd_sc_hd__xnor2_1 _12717_ (.A(_03533_),
    .B(_03534_),
    .Y(_03535_));
 sky130_fd_sc_hd__a32o_1 _12718_ (.A1(net417),
    .A2(net725),
    .A3(_03364_),
    .B1(_03365_),
    .B2(_03025_),
    .X(_03536_));
 sky130_fd_sc_hd__and2_2 _12719_ (.A(_03535_),
    .B(_03536_),
    .X(_03537_));
 sky130_fd_sc_hd__xor2_1 _12720_ (.A(_03535_),
    .B(_03536_),
    .X(_03539_));
 sky130_fd_sc_hd__a22oi_4 _12721_ (.A1(net442),
    .A2(net689),
    .B1(net699),
    .B2(net432),
    .Y(_03540_));
 sky130_fd_sc_hd__and4_1 _12722_ (.A(net432),
    .B(net442),
    .C(net689),
    .D(net699),
    .X(_03541_));
 sky130_fd_sc_hd__nor2_1 _12723_ (.A(_03540_),
    .B(_03541_),
    .Y(_03542_));
 sky130_fd_sc_hd__nand2_1 _12724_ (.A(net453),
    .B(net684),
    .Y(_03543_));
 sky130_fd_sc_hd__xnor2_1 _12725_ (.A(_03542_),
    .B(_03543_),
    .Y(_03544_));
 sky130_fd_sc_hd__and2_2 _12726_ (.A(_03539_),
    .B(_03544_),
    .X(_03545_));
 sky130_fd_sc_hd__nor2_1 _12727_ (.A(_03539_),
    .B(_03544_),
    .Y(_03546_));
 sky130_fd_sc_hd__or2_2 _12728_ (.A(_03545_),
    .B(_03546_),
    .X(_03547_));
 sky130_fd_sc_hd__a21o_4 _12729_ (.A1(_03370_),
    .A2(_03377_),
    .B1(_03547_),
    .X(_03548_));
 sky130_fd_sc_hd__nand3_2 _12730_ (.A(_03370_),
    .B(_03377_),
    .C(_03547_),
    .Y(_03550_));
 sky130_fd_sc_hd__o21ba_4 _12731_ (.A1(_03383_),
    .A2(_03386_),
    .B1_N(_03384_),
    .X(_03551_));
 sky130_fd_sc_hd__o21ba_4 _12732_ (.A1(_03372_),
    .A2(_03375_),
    .B1_N(_03373_),
    .X(_03552_));
 sky130_fd_sc_hd__a22oi_4 _12733_ (.A1(net469),
    .A2(net663),
    .B1(net671),
    .B2(net460),
    .Y(_03553_));
 sky130_fd_sc_hd__and4_1 _12734_ (.A(net460),
    .B(net469),
    .C(net663),
    .D(net671),
    .X(_03554_));
 sky130_fd_sc_hd__nor2_2 _12735_ (.A(_03553_),
    .B(_03554_),
    .Y(_03555_));
 sky130_fd_sc_hd__nand2_4 _12736_ (.A(net479),
    .B(net655),
    .Y(_03556_));
 sky130_fd_sc_hd__xnor2_4 _12737_ (.A(_03555_),
    .B(_03556_),
    .Y(_03557_));
 sky130_fd_sc_hd__and2b_1 _12738_ (.A_N(_03552_),
    .B(_03557_),
    .X(_03558_));
 sky130_fd_sc_hd__xnor2_4 _12739_ (.A(_03552_),
    .B(_03557_),
    .Y(_03559_));
 sky130_fd_sc_hd__and2b_1 _12740_ (.A_N(_03551_),
    .B(_03559_),
    .X(_03561_));
 sky130_fd_sc_hd__xnor2_4 _12741_ (.A(_03551_),
    .B(_03559_),
    .Y(_03562_));
 sky130_fd_sc_hd__a21o_1 _12742_ (.A1(_03548_),
    .A2(_03550_),
    .B1(_03562_),
    .X(_03563_));
 sky130_fd_sc_hd__nand3_4 _12743_ (.A(_03548_),
    .B(_03550_),
    .C(_03562_),
    .Y(_03564_));
 sky130_fd_sc_hd__and2_4 _12744_ (.A(_03563_),
    .B(_03564_),
    .X(_03565_));
 sky130_fd_sc_hd__a21bo_4 _12745_ (.A1(_03380_),
    .A2(_03392_),
    .B1_N(_03379_),
    .X(_03566_));
 sky130_fd_sc_hd__nand2_2 _12746_ (.A(_03565_),
    .B(_03566_),
    .Y(_03567_));
 sky130_fd_sc_hd__xnor2_4 _12747_ (.A(_03565_),
    .B(_03566_),
    .Y(_03568_));
 sky130_fd_sc_hd__a22oi_1 _12748_ (.A1(net494),
    .A2(net635),
    .B1(net645),
    .B2(net484),
    .Y(_03569_));
 sky130_fd_sc_hd__nand2_1 _12749_ (.A(net484),
    .B(net635),
    .Y(_03570_));
 sky130_fd_sc_hd__and4_2 _12750_ (.A(net485),
    .B(net494),
    .C(net635),
    .D(net645),
    .X(_03572_));
 sky130_fd_sc_hd__nor2_1 _12751_ (.A(_03569_),
    .B(_03572_),
    .Y(_03573_));
 sky130_fd_sc_hd__nand2_1 _12752_ (.A(net503),
    .B(net627),
    .Y(_03574_));
 sky130_fd_sc_hd__and3_2 _12753_ (.A(net503),
    .B(net627),
    .C(_03573_),
    .X(_03575_));
 sky130_fd_sc_hd__xnor2_1 _12754_ (.A(_03573_),
    .B(_03574_),
    .Y(_03576_));
 sky130_fd_sc_hd__or3_1 _12755_ (.A(_03405_),
    .B(_03409_),
    .C(_03576_),
    .X(_03577_));
 sky130_fd_sc_hd__o21ai_2 _12756_ (.A1(_03405_),
    .A2(_03409_),
    .B1(_03576_),
    .Y(_03578_));
 sky130_fd_sc_hd__and2_1 _12757_ (.A(_03577_),
    .B(_03578_),
    .X(_03579_));
 sky130_fd_sc_hd__nand2b_1 _12758_ (.A_N(_03401_),
    .B(_03579_),
    .Y(_03580_));
 sky130_fd_sc_hd__xnor2_1 _12759_ (.A(_03401_),
    .B(_03579_),
    .Y(_03581_));
 sky130_fd_sc_hd__o21a_1 _12760_ (.A1(_03389_),
    .A2(_03391_),
    .B1(_03581_),
    .X(_03583_));
 sky130_fd_sc_hd__nor3_1 _12761_ (.A(_03389_),
    .B(_03391_),
    .C(_03581_),
    .Y(_03584_));
 sky130_fd_sc_hd__or2_2 _12762_ (.A(_03583_),
    .B(_03584_),
    .X(_03585_));
 sky130_fd_sc_hd__a21oi_4 _12763_ (.A1(_03412_),
    .A2(_03414_),
    .B1(_03585_),
    .Y(_03586_));
 sky130_fd_sc_hd__and3_2 _12764_ (.A(_03412_),
    .B(_03414_),
    .C(_03585_),
    .X(_03587_));
 sky130_fd_sc_hd__o21ai_4 _12765_ (.A1(_03586_),
    .A2(_03587_),
    .B1(_03568_),
    .Y(_03588_));
 sky130_fd_sc_hd__or3_4 _12766_ (.A(_03568_),
    .B(_03586_),
    .C(_03587_),
    .X(_03589_));
 sky130_fd_sc_hd__o211ai_4 _12767_ (.A1(_03396_),
    .A2(_03423_),
    .B1(_03588_),
    .C1(_03589_),
    .Y(_03590_));
 sky130_fd_sc_hd__a211o_2 _12768_ (.A1(_03588_),
    .A2(_03589_),
    .B1(_03396_),
    .C1(_03423_),
    .X(_03591_));
 sky130_fd_sc_hd__a22oi_2 _12769_ (.A1(net328),
    .A2(net823),
    .B1(net831),
    .B2(net318),
    .Y(_03592_));
 sky130_fd_sc_hd__and4_1 _12770_ (.A(net318),
    .B(net328),
    .C(net823),
    .D(net831),
    .X(_03594_));
 sky130_fd_sc_hd__nor2_1 _12771_ (.A(_03592_),
    .B(_03594_),
    .Y(_03595_));
 sky130_fd_sc_hd__nand2_1 _12772_ (.A(net337),
    .B(net812),
    .Y(_03596_));
 sky130_fd_sc_hd__xnor2_1 _12773_ (.A(_03595_),
    .B(_03596_),
    .Y(_03597_));
 sky130_fd_sc_hd__and2_1 _12774_ (.A(_03402_),
    .B(_03597_),
    .X(_03598_));
 sky130_fd_sc_hd__nor2_1 _12775_ (.A(_03402_),
    .B(_03597_),
    .Y(_03599_));
 sky130_fd_sc_hd__or2_1 _12776_ (.A(_03598_),
    .B(_03599_),
    .X(_03600_));
 sky130_fd_sc_hd__a21oi_1 _12777_ (.A1(_03416_),
    .A2(_03419_),
    .B1(_03600_),
    .Y(_03601_));
 sky130_fd_sc_hd__and3_1 _12778_ (.A(_03416_),
    .B(_03419_),
    .C(_03600_),
    .X(_03602_));
 sky130_fd_sc_hd__nor2_2 _12779_ (.A(_03601_),
    .B(_03602_),
    .Y(_03603_));
 sky130_fd_sc_hd__xnor2_4 _12780_ (.A(_03434_),
    .B(_03603_),
    .Y(_03605_));
 sky130_fd_sc_hd__a21o_2 _12781_ (.A1(_03590_),
    .A2(_03591_),
    .B1(_03605_),
    .X(_03606_));
 sky130_fd_sc_hd__nand3_4 _12782_ (.A(_03590_),
    .B(_03591_),
    .C(_03605_),
    .Y(_03607_));
 sky130_fd_sc_hd__o211a_4 _12783_ (.A1(_03424_),
    .A2(_03443_),
    .B1(_03606_),
    .C1(_03607_),
    .X(_03608_));
 sky130_fd_sc_hd__a211oi_4 _12784_ (.A1(_03606_),
    .A2(_03607_),
    .B1(_03424_),
    .C1(_03443_),
    .Y(_03609_));
 sky130_fd_sc_hd__a32o_2 _12785_ (.A1(_03467_),
    .A2(_03468_),
    .A3(_03485_),
    .B1(_03483_),
    .B2(_03317_),
    .X(_03610_));
 sky130_fd_sc_hd__a22oi_4 _12786_ (.A1(net376),
    .A2(net761),
    .B1(net773),
    .B2(net367),
    .Y(_03611_));
 sky130_fd_sc_hd__and4_2 _12787_ (.A(net367),
    .B(net376),
    .C(net761),
    .D(net773),
    .X(_03612_));
 sky130_fd_sc_hd__nand2_1 _12788_ (.A(net384),
    .B(net751),
    .Y(_03613_));
 sky130_fd_sc_hd__o21a_1 _12789_ (.A1(_03611_),
    .A2(_03612_),
    .B1(_03613_),
    .X(_03614_));
 sky130_fd_sc_hd__nor3_2 _12790_ (.A(_03611_),
    .B(_03612_),
    .C(_03613_),
    .Y(_03616_));
 sky130_fd_sc_hd__nor2_2 _12791_ (.A(_03614_),
    .B(_03616_),
    .Y(_03617_));
 sky130_fd_sc_hd__nor3_2 _12792_ (.A(_03449_),
    .B(_03453_),
    .C(_03617_),
    .Y(_03618_));
 sky130_fd_sc_hd__o21a_2 _12793_ (.A1(_03449_),
    .A2(_03453_),
    .B1(_03617_),
    .X(_03619_));
 sky130_fd_sc_hd__nor2_4 _12794_ (.A(_03618_),
    .B(_03619_),
    .Y(_03620_));
 sky130_fd_sc_hd__nand2_2 _12795_ (.A(net389),
    .B(net738),
    .Y(_03621_));
 sky130_fd_sc_hd__xor2_4 _12796_ (.A(_03620_),
    .B(_03621_),
    .X(_03622_));
 sky130_fd_sc_hd__a21oi_4 _12797_ (.A1(_03456_),
    .A2(_03458_),
    .B1(_03622_),
    .Y(_03623_));
 sky130_fd_sc_hd__and3_1 _12798_ (.A(_03456_),
    .B(_03458_),
    .C(_03622_),
    .X(_03624_));
 sky130_fd_sc_hd__nor2_4 _12799_ (.A(_03623_),
    .B(_03624_),
    .Y(_03625_));
 sky130_fd_sc_hd__nand2_2 _12800_ (.A(net399),
    .B(net730),
    .Y(_03627_));
 sky130_fd_sc_hd__xnor2_4 _12801_ (.A(_03625_),
    .B(_03627_),
    .Y(_03628_));
 sky130_fd_sc_hd__o21ba_4 _12802_ (.A1(_03428_),
    .A2(_03432_),
    .B1_N(_03429_),
    .X(_03629_));
 sky130_fd_sc_hd__a22oi_4 _12803_ (.A1(net352),
    .A2(net795),
    .B1(net802),
    .B2(net344),
    .Y(_03630_));
 sky130_fd_sc_hd__and4_1 _12804_ (.A(net344),
    .B(net352),
    .C(net795),
    .D(net802),
    .X(_03631_));
 sky130_fd_sc_hd__nor2_2 _12805_ (.A(_03630_),
    .B(_03631_),
    .Y(_03632_));
 sky130_fd_sc_hd__nand2_4 _12806_ (.A(net359),
    .B(net779),
    .Y(_03633_));
 sky130_fd_sc_hd__xnor2_4 _12807_ (.A(_03632_),
    .B(_03633_),
    .Y(_03634_));
 sky130_fd_sc_hd__and2b_1 _12808_ (.A_N(_03629_),
    .B(_03634_),
    .X(_03635_));
 sky130_fd_sc_hd__xnor2_4 _12809_ (.A(_03629_),
    .B(_03634_),
    .Y(_03636_));
 sky130_fd_sc_hd__o21ba_2 _12810_ (.A1(_03470_),
    .A2(_03473_),
    .B1_N(_03471_),
    .X(_03638_));
 sky130_fd_sc_hd__and2b_1 _12811_ (.A_N(_03638_),
    .B(_03636_),
    .X(_03639_));
 sky130_fd_sc_hd__xor2_4 _12812_ (.A(_03636_),
    .B(_03638_),
    .X(_03640_));
 sky130_fd_sc_hd__o21ba_4 _12813_ (.A1(_03476_),
    .A2(_03478_),
    .B1_N(_03475_),
    .X(_03641_));
 sky130_fd_sc_hd__xor2_4 _12814_ (.A(_03640_),
    .B(_03641_),
    .X(_03642_));
 sky130_fd_sc_hd__nand2b_1 _12815_ (.A_N(_03481_),
    .B(_03642_),
    .Y(_03643_));
 sky130_fd_sc_hd__xnor2_2 _12816_ (.A(_03481_),
    .B(_03642_),
    .Y(_03644_));
 sky130_fd_sc_hd__xnor2_2 _12817_ (.A(_03628_),
    .B(_03644_),
    .Y(_03645_));
 sky130_fd_sc_hd__a21oi_1 _12818_ (.A1(_03437_),
    .A2(_03440_),
    .B1(_03645_),
    .Y(_03646_));
 sky130_fd_sc_hd__a21o_1 _12819_ (.A1(_03437_),
    .A2(_03440_),
    .B1(_03645_),
    .X(_03647_));
 sky130_fd_sc_hd__and3_1 _12820_ (.A(_03437_),
    .B(_03440_),
    .C(_03645_),
    .X(_03649_));
 sky130_fd_sc_hd__or2_1 _12821_ (.A(_03646_),
    .B(_03649_),
    .X(_03650_));
 sky130_fd_sc_hd__nand2b_4 _12822_ (.A_N(_03650_),
    .B(_03610_),
    .Y(_03651_));
 sky130_fd_sc_hd__nand2b_1 _12823_ (.A_N(_03610_),
    .B(_03650_),
    .Y(_03652_));
 sky130_fd_sc_hd__nand2_2 _12824_ (.A(_03651_),
    .B(_03652_),
    .Y(_03653_));
 sky130_fd_sc_hd__or3_4 _12825_ (.A(_03608_),
    .B(_03609_),
    .C(_03653_),
    .X(_03654_));
 sky130_fd_sc_hd__clkinv_2 _12826_ (.A(_03654_),
    .Y(_03655_));
 sky130_fd_sc_hd__o21ai_4 _12827_ (.A1(_03608_),
    .A2(_03609_),
    .B1(_03653_),
    .Y(_03656_));
 sky130_fd_sc_hd__o211a_2 _12828_ (.A1(_03444_),
    .A2(_03492_),
    .B1(_03654_),
    .C1(_03656_),
    .X(_03657_));
 sky130_fd_sc_hd__a211oi_4 _12829_ (.A1(_03654_),
    .A2(_03656_),
    .B1(_03444_),
    .C1(_03492_),
    .Y(_03658_));
 sky130_fd_sc_hd__a211oi_4 _12830_ (.A1(_03487_),
    .A2(_03489_),
    .B1(_03657_),
    .C1(_03658_),
    .Y(_03660_));
 sky130_fd_sc_hd__o211a_2 _12831_ (.A1(_03657_),
    .A2(_03658_),
    .B1(_03487_),
    .C1(_03489_),
    .X(_03661_));
 sky130_fd_sc_hd__o21ba_2 _12832_ (.A1(_03498_),
    .A2(_03499_),
    .B1_N(_03497_),
    .X(_03662_));
 sky130_fd_sc_hd__nor3_4 _12833_ (.A(_03660_),
    .B(_03661_),
    .C(_03662_),
    .Y(_03663_));
 sky130_fd_sc_hd__or3_4 _12834_ (.A(_03660_),
    .B(_03661_),
    .C(_03662_),
    .X(_03664_));
 sky130_fd_sc_hd__o21a_2 _12835_ (.A1(_03660_),
    .A2(_03661_),
    .B1(_03662_),
    .X(_03665_));
 sky130_fd_sc_hd__a211o_4 _12836_ (.A1(_03462_),
    .A2(_03467_),
    .B1(_03663_),
    .C1(_03665_),
    .X(_03666_));
 sky130_fd_sc_hd__o211ai_4 _12837_ (.A1(_03663_),
    .A2(_03665_),
    .B1(_03462_),
    .C1(_03467_),
    .Y(_03667_));
 sky130_fd_sc_hd__a211oi_4 _12838_ (.A1(_03666_),
    .A2(_03667_),
    .B1(_03502_),
    .C1(_03505_),
    .Y(_03668_));
 sky130_fd_sc_hd__o211ai_4 _12839_ (.A1(_03502_),
    .A2(_03505_),
    .B1(_03666_),
    .C1(_03667_),
    .Y(_03669_));
 sky130_fd_sc_hd__nand2b_2 _12840_ (.A_N(_03668_),
    .B(_03669_),
    .Y(_03671_));
 sky130_fd_sc_hd__o21ai_1 _12841_ (.A1(_03511_),
    .A2(_03514_),
    .B1(_03510_),
    .Y(_03672_));
 sky130_fd_sc_hd__xnor2_1 _12842_ (.A(_03671_),
    .B(_03672_),
    .Y(_03673_));
 sky130_fd_sc_hd__nand2_1 _12843_ (.A(net260),
    .B(_03673_),
    .Y(_03674_));
 sky130_fd_sc_hd__mux2_1 _12844_ (.A0(_03014_),
    .A1(_03016_),
    .S(net293),
    .X(_03675_));
 sky130_fd_sc_hd__mux2_2 _12845_ (.A0(_03004_),
    .A1(_03017_),
    .S(net584),
    .X(_03676_));
 sky130_fd_sc_hd__mux2_1 _12846_ (.A0(_03675_),
    .A1(_03676_),
    .S(net300),
    .X(_03677_));
 sky130_fd_sc_hd__and2_1 _12847_ (.A(net552),
    .B(_03677_),
    .X(_03678_));
 sky130_fd_sc_hd__mux2_2 _12848_ (.A0(_03005_),
    .A1(_03009_),
    .S(net293),
    .X(_03679_));
 sky130_fd_sc_hd__or2_1 _12849_ (.A(net300),
    .B(_03679_),
    .X(_03680_));
 sky130_fd_sc_hd__a211o_1 _12850_ (.A1(net305),
    .A2(_03680_),
    .B1(_03678_),
    .C1(net208),
    .X(_03682_));
 sky130_fd_sc_hd__mux2_1 _12851_ (.A0(_03013_),
    .A1(_03021_),
    .S(net584),
    .X(_03683_));
 sky130_fd_sc_hd__or2_4 _12852_ (.A(net570),
    .B(_03683_),
    .X(_03684_));
 sky130_fd_sc_hd__and2_2 _12853_ (.A(net538),
    .B(_02641_),
    .X(_03685_));
 sky130_fd_sc_hd__nand2_1 _12854_ (.A(net537),
    .B(_02641_),
    .Y(_03686_));
 sky130_fd_sc_hd__o31a_1 _12855_ (.A1(net563),
    .A2(_03684_),
    .A3(net205),
    .B1(_03682_),
    .X(_03687_));
 sky130_fd_sc_hd__nand2_1 _12856_ (.A(_03674_),
    .B(_03687_),
    .Y(_08680_));
 sky130_fd_sc_hd__mux2_1 _12857_ (.A0(_03174_),
    .A1(_03191_),
    .S(net585),
    .X(_03688_));
 sky130_fd_sc_hd__nand2_8 _12858_ (.A(net567),
    .B(net295),
    .Y(_03689_));
 sky130_fd_sc_hd__o22a_1 _12859_ (.A1(net568),
    .A2(_03688_),
    .B1(_03689_),
    .B2(_03190_),
    .X(_03690_));
 sky130_fd_sc_hd__o21ai_1 _12860_ (.A1(net206),
    .A2(_03690_),
    .B1(net209),
    .Y(_03692_));
 sky130_fd_sc_hd__mux2_1 _12861_ (.A0(_03175_),
    .A1(_03177_),
    .S(net296),
    .X(_03693_));
 sky130_fd_sc_hd__mux2_1 _12862_ (.A0(_03178_),
    .A1(_03181_),
    .S(net296),
    .X(_03694_));
 sky130_fd_sc_hd__mux2_1 _12863_ (.A0(_03693_),
    .A1(_03694_),
    .S(net301),
    .X(_03695_));
 sky130_fd_sc_hd__inv_2 _12864_ (.A(_03695_),
    .Y(_03696_));
 sky130_fd_sc_hd__mux2_1 _12865_ (.A0(_03183_),
    .A1(_03185_),
    .S(net295),
    .X(_03697_));
 sky130_fd_sc_hd__nor2_1 _12866_ (.A(net552),
    .B(_03697_),
    .Y(_03698_));
 sky130_fd_sc_hd__a221o_1 _12867_ (.A1(net552),
    .A2(_03696_),
    .B1(_03698_),
    .B2(net568),
    .C1(net537),
    .X(_03699_));
 sky130_fd_sc_hd__a21oi_2 _12868_ (.A1(net423),
    .A2(net699),
    .B1(_03365_),
    .Y(_03700_));
 sky130_fd_sc_hd__and3_2 _12869_ (.A(net423),
    .B(net699),
    .C(_03365_),
    .X(_03701_));
 sky130_fd_sc_hd__nor2_4 _12870_ (.A(_03700_),
    .B(_03701_),
    .Y(_03703_));
 sky130_fd_sc_hd__nand2_2 _12871_ (.A(net416),
    .B(net706),
    .Y(_03704_));
 sky130_fd_sc_hd__xnor2_4 _12872_ (.A(_03703_),
    .B(_03704_),
    .Y(_03705_));
 sky130_fd_sc_hd__o21ba_2 _12873_ (.A1(_03531_),
    .A2(_03534_),
    .B1_N(_03532_),
    .X(_03706_));
 sky130_fd_sc_hd__nand2b_2 _12874_ (.A_N(_03706_),
    .B(_03705_),
    .Y(_03707_));
 sky130_fd_sc_hd__xor2_4 _12875_ (.A(_03705_),
    .B(_03706_),
    .X(_03708_));
 sky130_fd_sc_hd__a22oi_1 _12876_ (.A1(net442),
    .A2(net684),
    .B1(net689),
    .B2(net432),
    .Y(_03709_));
 sky130_fd_sc_hd__and4_1 _12877_ (.A(net432),
    .B(net442),
    .C(net684),
    .D(net689),
    .X(_03710_));
 sky130_fd_sc_hd__or2_1 _12878_ (.A(_03709_),
    .B(_03710_),
    .X(_03711_));
 sky130_fd_sc_hd__nand2_1 _12879_ (.A(net453),
    .B(net671),
    .Y(_03712_));
 sky130_fd_sc_hd__nor2_1 _12880_ (.A(_03711_),
    .B(_03712_),
    .Y(_03714_));
 sky130_fd_sc_hd__nand2_1 _12881_ (.A(_03711_),
    .B(_03712_),
    .Y(_03715_));
 sky130_fd_sc_hd__and2b_4 _12882_ (.A_N(_03714_),
    .B(_03715_),
    .X(_03716_));
 sky130_fd_sc_hd__nand2b_2 _12883_ (.A_N(_03708_),
    .B(_03716_),
    .Y(_03717_));
 sky130_fd_sc_hd__xnor2_4 _12884_ (.A(_03708_),
    .B(_03716_),
    .Y(_03718_));
 sky130_fd_sc_hd__o21ai_4 _12885_ (.A1(_03537_),
    .A2(_03545_),
    .B1(_03718_),
    .Y(_03719_));
 sky130_fd_sc_hd__or3_4 _12886_ (.A(_03537_),
    .B(_03545_),
    .C(_03718_),
    .X(_03720_));
 sky130_fd_sc_hd__o21ba_2 _12887_ (.A1(_03553_),
    .A2(_03556_),
    .B1_N(_03554_),
    .X(_03721_));
 sky130_fd_sc_hd__o21ba_4 _12888_ (.A1(_03540_),
    .A2(_03543_),
    .B1_N(_03541_),
    .X(_03722_));
 sky130_fd_sc_hd__a22oi_2 _12889_ (.A1(net470),
    .A2(net654),
    .B1(net662),
    .B2(net459),
    .Y(_03723_));
 sky130_fd_sc_hd__and4_1 _12890_ (.A(net459),
    .B(net469),
    .C(net654),
    .D(net662),
    .X(_03725_));
 sky130_fd_sc_hd__and4bb_2 _12891_ (.A_N(_03723_),
    .B_N(_03725_),
    .C(net479),
    .D(net644),
    .X(_03726_));
 sky130_fd_sc_hd__o2bb2a_1 _12892_ (.A1_N(net479),
    .A2_N(net644),
    .B1(_03723_),
    .B2(_03725_),
    .X(_03727_));
 sky130_fd_sc_hd__nor2_4 _12893_ (.A(_03726_),
    .B(_03727_),
    .Y(_03728_));
 sky130_fd_sc_hd__and2b_1 _12894_ (.A_N(_03722_),
    .B(_03728_),
    .X(_03729_));
 sky130_fd_sc_hd__xnor2_4 _12895_ (.A(_03722_),
    .B(_03728_),
    .Y(_03730_));
 sky130_fd_sc_hd__and2b_1 _12896_ (.A_N(_03721_),
    .B(_03730_),
    .X(_03731_));
 sky130_fd_sc_hd__xnor2_4 _12897_ (.A(_03721_),
    .B(_03730_),
    .Y(_03732_));
 sky130_fd_sc_hd__a21o_1 _12898_ (.A1(_03719_),
    .A2(_03720_),
    .B1(_03732_),
    .X(_03733_));
 sky130_fd_sc_hd__nand3_4 _12899_ (.A(_03719_),
    .B(_03720_),
    .C(_03732_),
    .Y(_03734_));
 sky130_fd_sc_hd__nand2_2 _12900_ (.A(_03733_),
    .B(_03734_),
    .Y(_03736_));
 sky130_fd_sc_hd__a21o_4 _12901_ (.A1(_03548_),
    .A2(_03564_),
    .B1(_03736_),
    .X(_03737_));
 sky130_fd_sc_hd__nand3_4 _12902_ (.A(_03548_),
    .B(_03564_),
    .C(_03736_),
    .Y(_03738_));
 sky130_fd_sc_hd__or2_2 _12903_ (.A(_03558_),
    .B(_03561_),
    .X(_03739_));
 sky130_fd_sc_hd__nand2_2 _12904_ (.A(net495),
    .B(net627),
    .Y(_03740_));
 sky130_fd_sc_hd__and4_4 _12905_ (.A(net485),
    .B(net495),
    .C(net627),
    .D(net635),
    .X(_03741_));
 sky130_fd_sc_hd__a21oi_4 _12906_ (.A1(_03570_),
    .A2(_03740_),
    .B1(_03741_),
    .Y(_03742_));
 sky130_fd_sc_hd__nand2_1 _12907_ (.A(net503),
    .B(net619),
    .Y(_03743_));
 sky130_fd_sc_hd__xnor2_2 _12908_ (.A(_03742_),
    .B(_03743_),
    .Y(_03744_));
 sky130_fd_sc_hd__o21ai_4 _12909_ (.A1(_03572_),
    .A2(_03575_),
    .B1(_03744_),
    .Y(_03745_));
 sky130_fd_sc_hd__or3_1 _12910_ (.A(_03572_),
    .B(_03575_),
    .C(_03744_),
    .X(_03747_));
 sky130_fd_sc_hd__and2_1 _12911_ (.A(_03745_),
    .B(_03747_),
    .X(_03748_));
 sky130_fd_sc_hd__and2_1 _12912_ (.A(_03739_),
    .B(_03748_),
    .X(_03749_));
 sky130_fd_sc_hd__xnor2_1 _12913_ (.A(_03739_),
    .B(_03748_),
    .Y(_03750_));
 sky130_fd_sc_hd__a21oi_2 _12914_ (.A1(_03578_),
    .A2(_03580_),
    .B1(_03750_),
    .Y(_03751_));
 sky130_fd_sc_hd__and3_1 _12915_ (.A(_03578_),
    .B(_03580_),
    .C(_03750_),
    .X(_03752_));
 sky130_fd_sc_hd__nor2_2 _12916_ (.A(_03751_),
    .B(_03752_),
    .Y(_03753_));
 sky130_fd_sc_hd__a21o_1 _12917_ (.A1(_03737_),
    .A2(_03738_),
    .B1(_03753_),
    .X(_03754_));
 sky130_fd_sc_hd__nand3_4 _12918_ (.A(_03737_),
    .B(_03738_),
    .C(_03753_),
    .Y(_03755_));
 sky130_fd_sc_hd__nand2_2 _12919_ (.A(_03754_),
    .B(_03755_),
    .Y(_03756_));
 sky130_fd_sc_hd__and3_2 _12920_ (.A(_03567_),
    .B(_03589_),
    .C(_03756_),
    .X(_03758_));
 sky130_fd_sc_hd__a21oi_4 _12921_ (.A1(_03567_),
    .A2(_03589_),
    .B1(_03756_),
    .Y(_03759_));
 sky130_fd_sc_hd__a22oi_2 _12922_ (.A1(net328),
    .A2(net812),
    .B1(net823),
    .B2(net318),
    .Y(_03760_));
 sky130_fd_sc_hd__and4_1 _12923_ (.A(net318),
    .B(net328),
    .C(net812),
    .D(net823),
    .X(_03761_));
 sky130_fd_sc_hd__nor2_1 _12924_ (.A(_03760_),
    .B(_03761_),
    .Y(_03762_));
 sky130_fd_sc_hd__nand2_2 _12925_ (.A(net337),
    .B(net802),
    .Y(_03763_));
 sky130_fd_sc_hd__xnor2_2 _12926_ (.A(_03762_),
    .B(_03763_),
    .Y(_03764_));
 sky130_fd_sc_hd__o21ai_2 _12927_ (.A1(_03583_),
    .A2(_03586_),
    .B1(_03764_),
    .Y(_03765_));
 sky130_fd_sc_hd__or3_1 _12928_ (.A(_03583_),
    .B(_03586_),
    .C(_03764_),
    .X(_03766_));
 sky130_fd_sc_hd__and2_1 _12929_ (.A(_03765_),
    .B(_03766_),
    .X(_03767_));
 sky130_fd_sc_hd__nand2_2 _12930_ (.A(_03598_),
    .B(_03767_),
    .Y(_03769_));
 sky130_fd_sc_hd__or2_1 _12931_ (.A(_03598_),
    .B(_03767_),
    .X(_03770_));
 sky130_fd_sc_hd__nand2_2 _12932_ (.A(_03769_),
    .B(_03770_),
    .Y(_03771_));
 sky130_fd_sc_hd__nor3_4 _12933_ (.A(_03758_),
    .B(_03759_),
    .C(_03771_),
    .Y(_03772_));
 sky130_fd_sc_hd__o21a_1 _12934_ (.A1(_03758_),
    .A2(_03759_),
    .B1(_03771_),
    .X(_03773_));
 sky130_fd_sc_hd__or2_4 _12935_ (.A(_03772_),
    .B(_03773_),
    .X(_03774_));
 sky130_fd_sc_hd__a21oi_4 _12936_ (.A1(_03590_),
    .A2(_03607_),
    .B1(_03774_),
    .Y(_03775_));
 sky130_fd_sc_hd__inv_2 _12937_ (.A(_03775_),
    .Y(_03776_));
 sky130_fd_sc_hd__and3_2 _12938_ (.A(_03590_),
    .B(_03607_),
    .C(_03774_),
    .X(_03777_));
 sky130_fd_sc_hd__a21bo_2 _12939_ (.A1(_03628_),
    .A2(_03644_),
    .B1_N(_03643_),
    .X(_03778_));
 sky130_fd_sc_hd__o21ba_1 _12940_ (.A1(_03434_),
    .A2(_03602_),
    .B1_N(_03601_),
    .X(_03780_));
 sky130_fd_sc_hd__a22oi_4 _12941_ (.A1(net376),
    .A2(net751),
    .B1(net761),
    .B2(net367),
    .Y(_03781_));
 sky130_fd_sc_hd__and4_2 _12942_ (.A(net367),
    .B(net376),
    .C(net751),
    .D(net761),
    .X(_03782_));
 sky130_fd_sc_hd__nand2_1 _12943_ (.A(net384),
    .B(net742),
    .Y(_03783_));
 sky130_fd_sc_hd__o21a_1 _12944_ (.A1(_03781_),
    .A2(_03782_),
    .B1(_03783_),
    .X(_03784_));
 sky130_fd_sc_hd__nor3_2 _12945_ (.A(_03781_),
    .B(_03782_),
    .C(_03783_),
    .Y(_03785_));
 sky130_fd_sc_hd__nor2_1 _12946_ (.A(_03784_),
    .B(_03785_),
    .Y(_03786_));
 sky130_fd_sc_hd__or3_1 _12947_ (.A(_03612_),
    .B(_03616_),
    .C(_03786_),
    .X(_03787_));
 sky130_fd_sc_hd__o21ai_1 _12948_ (.A1(_03612_),
    .A2(_03616_),
    .B1(_03786_),
    .Y(_03788_));
 sky130_fd_sc_hd__and2_1 _12949_ (.A(_03787_),
    .B(_03788_),
    .X(_03789_));
 sky130_fd_sc_hd__nand3_1 _12950_ (.A(net393),
    .B(net733),
    .C(_03789_),
    .Y(_03791_));
 sky130_fd_sc_hd__a21o_1 _12951_ (.A1(net393),
    .A2(net733),
    .B1(_03789_),
    .X(_03792_));
 sky130_fd_sc_hd__nand2_1 _12952_ (.A(_03791_),
    .B(_03792_),
    .Y(_03793_));
 sky130_fd_sc_hd__a31o_1 _12953_ (.A1(net393),
    .A2(net738),
    .A3(_03620_),
    .B1(_03619_),
    .X(_03794_));
 sky130_fd_sc_hd__nand2b_2 _12954_ (.A_N(_03793_),
    .B(_03794_),
    .Y(_03795_));
 sky130_fd_sc_hd__nand2b_1 _12955_ (.A_N(_03794_),
    .B(_03793_),
    .Y(_03796_));
 sky130_fd_sc_hd__nand2_1 _12956_ (.A(_03795_),
    .B(_03796_),
    .Y(_03797_));
 sky130_fd_sc_hd__nand2_1 _12957_ (.A(net401),
    .B(net721),
    .Y(_03798_));
 sky130_fd_sc_hd__or2_2 _12958_ (.A(_03797_),
    .B(_03798_),
    .X(_03799_));
 sky130_fd_sc_hd__nand2_1 _12959_ (.A(_03797_),
    .B(_03798_),
    .Y(_03800_));
 sky130_fd_sc_hd__and2_2 _12960_ (.A(_03799_),
    .B(_03800_),
    .X(_03802_));
 sky130_fd_sc_hd__o21ba_1 _12961_ (.A1(_03592_),
    .A2(_03596_),
    .B1_N(_03594_),
    .X(_03803_));
 sky130_fd_sc_hd__a22oi_2 _12962_ (.A1(net352),
    .A2(net779),
    .B1(net795),
    .B2(net344),
    .Y(_03804_));
 sky130_fd_sc_hd__and4_1 _12963_ (.A(net344),
    .B(net352),
    .C(net779),
    .D(net795),
    .X(_03805_));
 sky130_fd_sc_hd__nor2_1 _12964_ (.A(_03804_),
    .B(_03805_),
    .Y(_03806_));
 sky130_fd_sc_hd__nand2_2 _12965_ (.A(net359),
    .B(net773),
    .Y(_03807_));
 sky130_fd_sc_hd__xnor2_2 _12966_ (.A(_03806_),
    .B(_03807_),
    .Y(_03808_));
 sky130_fd_sc_hd__and2b_1 _12967_ (.A_N(_03803_),
    .B(_03808_),
    .X(_03809_));
 sky130_fd_sc_hd__xnor2_1 _12968_ (.A(_03803_),
    .B(_03808_),
    .Y(_03810_));
 sky130_fd_sc_hd__o21ba_1 _12969_ (.A1(_03630_),
    .A2(_03633_),
    .B1_N(_03631_),
    .X(_03811_));
 sky130_fd_sc_hd__and2b_1 _12970_ (.A_N(_03811_),
    .B(_03810_),
    .X(_03813_));
 sky130_fd_sc_hd__xor2_1 _12971_ (.A(_03810_),
    .B(_03811_),
    .X(_03814_));
 sky130_fd_sc_hd__nor2_1 _12972_ (.A(_03635_),
    .B(_03639_),
    .Y(_03815_));
 sky130_fd_sc_hd__or2_2 _12973_ (.A(_03814_),
    .B(_03815_),
    .X(_03816_));
 sky130_fd_sc_hd__nand2_1 _12974_ (.A(_03814_),
    .B(_03815_),
    .Y(_03817_));
 sky130_fd_sc_hd__and2_1 _12975_ (.A(_03816_),
    .B(_03817_),
    .X(_03818_));
 sky130_fd_sc_hd__or3b_1 _12976_ (.A(_03640_),
    .B(_03641_),
    .C_N(_03818_),
    .X(_03819_));
 sky130_fd_sc_hd__o21bai_1 _12977_ (.A1(_03640_),
    .A2(_03641_),
    .B1_N(_03818_),
    .Y(_03820_));
 sky130_fd_sc_hd__and2_1 _12978_ (.A(_03819_),
    .B(_03820_),
    .X(_03821_));
 sky130_fd_sc_hd__xnor2_2 _12979_ (.A(_03802_),
    .B(_03821_),
    .Y(_03822_));
 sky130_fd_sc_hd__or2_4 _12980_ (.A(_03780_),
    .B(_03822_),
    .X(_03824_));
 sky130_fd_sc_hd__xnor2_1 _12981_ (.A(_03780_),
    .B(_03822_),
    .Y(_03825_));
 sky130_fd_sc_hd__nand2b_4 _12982_ (.A_N(_03825_),
    .B(_03778_),
    .Y(_03826_));
 sky130_fd_sc_hd__nand2b_1 _12983_ (.A_N(_03778_),
    .B(_03825_),
    .Y(_03827_));
 sky130_fd_sc_hd__nand2_2 _12984_ (.A(_03826_),
    .B(_03827_),
    .Y(_03828_));
 sky130_fd_sc_hd__or3_4 _12985_ (.A(_03775_),
    .B(_03777_),
    .C(_03828_),
    .X(_03829_));
 sky130_fd_sc_hd__o21ai_4 _12986_ (.A1(_03775_),
    .A2(_03777_),
    .B1(_03828_),
    .Y(_03830_));
 sky130_fd_sc_hd__o211a_4 _12987_ (.A1(_03608_),
    .A2(_03655_),
    .B1(_03829_),
    .C1(_03830_),
    .X(_03831_));
 sky130_fd_sc_hd__a211oi_4 _12988_ (.A1(_03829_),
    .A2(_03830_),
    .B1(_03608_),
    .C1(_03655_),
    .Y(_03832_));
 sky130_fd_sc_hd__a211oi_4 _12989_ (.A1(_03647_),
    .A2(_03651_),
    .B1(_03831_),
    .C1(_03832_),
    .Y(_03833_));
 sky130_fd_sc_hd__o211a_1 _12990_ (.A1(_03831_),
    .A2(_03832_),
    .B1(_03647_),
    .C1(_03651_),
    .X(_03835_));
 sky130_fd_sc_hd__or2_1 _12991_ (.A(_03657_),
    .B(_03660_),
    .X(_03836_));
 sky130_fd_sc_hd__nor3b_1 _12992_ (.A(_03833_),
    .B(_03835_),
    .C_N(_03836_),
    .Y(_03837_));
 sky130_fd_sc_hd__or3b_1 _12993_ (.A(_03833_),
    .B(_03835_),
    .C_N(_03836_),
    .X(_03838_));
 sky130_fd_sc_hd__o21ba_1 _12994_ (.A1(_03833_),
    .A2(_03835_),
    .B1_N(_03836_),
    .X(_03839_));
 sky130_fd_sc_hd__a31o_1 _12995_ (.A1(net399),
    .A2(net730),
    .A3(_03625_),
    .B1(_03623_),
    .X(_03840_));
 sky130_fd_sc_hd__inv_2 _12996_ (.A(_03840_),
    .Y(_03841_));
 sky130_fd_sc_hd__or3_2 _12997_ (.A(_03837_),
    .B(_03839_),
    .C(_03841_),
    .X(_03842_));
 sky130_fd_sc_hd__o21ai_1 _12998_ (.A1(_03837_),
    .A2(_03839_),
    .B1(_03841_),
    .Y(_03843_));
 sky130_fd_sc_hd__nand2_2 _12999_ (.A(_03842_),
    .B(_03843_),
    .Y(_03844_));
 sky130_fd_sc_hd__a21oi_4 _13000_ (.A1(_03664_),
    .A2(_03666_),
    .B1(_03844_),
    .Y(_03846_));
 sky130_fd_sc_hd__and3_1 _13001_ (.A(_03664_),
    .B(_03666_),
    .C(_03844_),
    .X(_03847_));
 sky130_fd_sc_hd__or2_1 _13002_ (.A(_03846_),
    .B(_03847_),
    .X(_03848_));
 sky130_fd_sc_hd__or2_1 _13003_ (.A(_03511_),
    .B(_03671_),
    .X(_03849_));
 sky130_fd_sc_hd__nor2_1 _13004_ (.A(_03513_),
    .B(_03849_),
    .Y(_03850_));
 sky130_fd_sc_hd__and2_1 _13005_ (.A(_03168_),
    .B(_03850_),
    .X(_03851_));
 sky130_fd_sc_hd__a21oi_1 _13006_ (.A1(_03510_),
    .A2(_03669_),
    .B1(_03668_),
    .Y(_03852_));
 sky130_fd_sc_hd__o21bai_1 _13007_ (.A1(_03512_),
    .A2(_03849_),
    .B1_N(_03852_),
    .Y(_03853_));
 sky130_fd_sc_hd__a311o_4 _13008_ (.A1(_02574_),
    .A2(_03169_),
    .A3(_03850_),
    .B1(_03851_),
    .C1(_03853_),
    .X(_03854_));
 sky130_fd_sc_hd__nand2b_1 _13009_ (.A_N(_03854_),
    .B(_03848_),
    .Y(_03855_));
 sky130_fd_sc_hd__nand2b_1 _13010_ (.A_N(_03848_),
    .B(_03854_),
    .Y(_03857_));
 sky130_fd_sc_hd__a32o_1 _13011_ (.A1(net260),
    .A2(_03855_),
    .A3(_03857_),
    .B1(_03692_),
    .B2(_03699_),
    .X(_08681_));
 sky130_fd_sc_hd__o22a_4 _13012_ (.A1(net567),
    .A2(_02628_),
    .B1(_02647_),
    .B2(_03689_),
    .X(_03858_));
 sky130_fd_sc_hd__o21ai_1 _13013_ (.A1(net206),
    .A2(_03858_),
    .B1(net209),
    .Y(_03859_));
 sky130_fd_sc_hd__mux4_2 _13014_ (.A0(_02600_),
    .A1(_02605_),
    .A2(_02633_),
    .A3(_02638_),
    .S0(net293),
    .S1(net567),
    .X(_03860_));
 sky130_fd_sc_hd__nor2_1 _13015_ (.A(net307),
    .B(_03860_),
    .Y(_03861_));
 sky130_fd_sc_hd__a311o_1 _13016_ (.A1(net307),
    .A2(net570),
    .A3(_02614_),
    .B1(_03861_),
    .C1(net539),
    .X(_03862_));
 sky130_fd_sc_hd__a22oi_4 _13017_ (.A1(net423),
    .A2(net690),
    .B1(net707),
    .B2(net407),
    .Y(_03863_));
 sky130_fd_sc_hd__and4_1 _13018_ (.A(net407),
    .B(net423),
    .C(net690),
    .D(net707),
    .X(_03864_));
 sky130_fd_sc_hd__nor2_2 _13019_ (.A(_03863_),
    .B(_03864_),
    .Y(_03865_));
 sky130_fd_sc_hd__nand2_4 _13020_ (.A(net416),
    .B(net698),
    .Y(_03867_));
 sky130_fd_sc_hd__xnor2_4 _13021_ (.A(_03865_),
    .B(_03867_),
    .Y(_03868_));
 sky130_fd_sc_hd__a31o_4 _13022_ (.A1(net416),
    .A2(net706),
    .A3(_03703_),
    .B1(_03701_),
    .X(_03869_));
 sky130_fd_sc_hd__nand2_2 _13023_ (.A(_03868_),
    .B(_03869_),
    .Y(_03870_));
 sky130_fd_sc_hd__xor2_4 _13024_ (.A(_03868_),
    .B(_03869_),
    .X(_03871_));
 sky130_fd_sc_hd__a22oi_4 _13025_ (.A1(net442),
    .A2(net670),
    .B1(net680),
    .B2(net432),
    .Y(_03872_));
 sky130_fd_sc_hd__and4_1 _13026_ (.A(net432),
    .B(net442),
    .C(net670),
    .D(net680),
    .X(_03873_));
 sky130_fd_sc_hd__nor2_2 _13027_ (.A(_03872_),
    .B(_03873_),
    .Y(_03874_));
 sky130_fd_sc_hd__nand2_4 _13028_ (.A(net450),
    .B(net662),
    .Y(_03875_));
 sky130_fd_sc_hd__xnor2_4 _13029_ (.A(_03874_),
    .B(_03875_),
    .Y(_03876_));
 sky130_fd_sc_hd__nand2_2 _13030_ (.A(_03871_),
    .B(_03876_),
    .Y(_03878_));
 sky130_fd_sc_hd__xnor2_2 _13031_ (.A(_03871_),
    .B(_03876_),
    .Y(_03879_));
 sky130_fd_sc_hd__a21o_4 _13032_ (.A1(_03707_),
    .A2(_03717_),
    .B1(_03879_),
    .X(_03880_));
 sky130_fd_sc_hd__nand3_2 _13033_ (.A(_03707_),
    .B(_03717_),
    .C(_03879_),
    .Y(_03881_));
 sky130_fd_sc_hd__a22oi_4 _13034_ (.A1(net470),
    .A2(net644),
    .B1(net654),
    .B2(net459),
    .Y(_03882_));
 sky130_fd_sc_hd__and4_1 _13035_ (.A(net459),
    .B(net470),
    .C(net644),
    .D(net654),
    .X(_03883_));
 sky130_fd_sc_hd__nor2_1 _13036_ (.A(_03882_),
    .B(_03883_),
    .Y(_03884_));
 sky130_fd_sc_hd__nand2_1 _13037_ (.A(net479),
    .B(net635),
    .Y(_03885_));
 sky130_fd_sc_hd__xnor2_1 _13038_ (.A(_03884_),
    .B(_03885_),
    .Y(_03886_));
 sky130_fd_sc_hd__o21ai_1 _13039_ (.A1(_03710_),
    .A2(_03714_),
    .B1(_03886_),
    .Y(_03887_));
 sky130_fd_sc_hd__or3_1 _13040_ (.A(_03710_),
    .B(_03714_),
    .C(_03886_),
    .X(_03889_));
 sky130_fd_sc_hd__and2_1 _13041_ (.A(_03887_),
    .B(_03889_),
    .X(_03890_));
 sky130_fd_sc_hd__o21ai_1 _13042_ (.A1(_03725_),
    .A2(_03726_),
    .B1(_03890_),
    .Y(_03891_));
 sky130_fd_sc_hd__or3_1 _13043_ (.A(_03725_),
    .B(_03726_),
    .C(_03890_),
    .X(_03892_));
 sky130_fd_sc_hd__and2_2 _13044_ (.A(_03891_),
    .B(_03892_),
    .X(_03893_));
 sky130_fd_sc_hd__a21o_1 _13045_ (.A1(_03880_),
    .A2(_03881_),
    .B1(_03893_),
    .X(_03894_));
 sky130_fd_sc_hd__nand3_4 _13046_ (.A(_03880_),
    .B(_03881_),
    .C(_03893_),
    .Y(_03895_));
 sky130_fd_sc_hd__nand2_1 _13047_ (.A(_03894_),
    .B(_03895_),
    .Y(_03896_));
 sky130_fd_sc_hd__a21o_4 _13048_ (.A1(_03719_),
    .A2(_03734_),
    .B1(_03896_),
    .X(_03897_));
 sky130_fd_sc_hd__nand3_2 _13049_ (.A(_03719_),
    .B(_03734_),
    .C(_03896_),
    .Y(_03898_));
 sky130_fd_sc_hd__a22oi_1 _13050_ (.A1(net495),
    .A2(net619),
    .B1(net627),
    .B2(net485),
    .Y(_03900_));
 sky130_fd_sc_hd__and4_2 _13051_ (.A(net485),
    .B(net495),
    .C(net619),
    .D(net627),
    .X(_03901_));
 sky130_fd_sc_hd__or2_2 _13052_ (.A(_03900_),
    .B(_03901_),
    .X(_03902_));
 sky130_fd_sc_hd__a31oi_4 _13053_ (.A1(net503),
    .A2(net619),
    .A3(_03742_),
    .B1(_03741_),
    .Y(_03903_));
 sky130_fd_sc_hd__or2_1 _13054_ (.A(_03902_),
    .B(_03903_),
    .X(_03904_));
 sky130_fd_sc_hd__xor2_2 _13055_ (.A(_03902_),
    .B(_03903_),
    .X(_03905_));
 sky130_fd_sc_hd__o21a_2 _13056_ (.A1(_03729_),
    .A2(_03731_),
    .B1(_03905_),
    .X(_03906_));
 sky130_fd_sc_hd__nor3_2 _13057_ (.A(_03729_),
    .B(_03731_),
    .C(_03905_),
    .Y(_03907_));
 sky130_fd_sc_hd__nor2_4 _13058_ (.A(_03906_),
    .B(_03907_),
    .Y(_03908_));
 sky130_fd_sc_hd__and2b_1 _13059_ (.A_N(_03745_),
    .B(_03908_),
    .X(_03909_));
 sky130_fd_sc_hd__xnor2_4 _13060_ (.A(_03745_),
    .B(_03908_),
    .Y(_03911_));
 sky130_fd_sc_hd__nand3_4 _13061_ (.A(_03897_),
    .B(_03898_),
    .C(_03911_),
    .Y(_03912_));
 sky130_fd_sc_hd__a21o_1 _13062_ (.A1(_03897_),
    .A2(_03898_),
    .B1(_03911_),
    .X(_03913_));
 sky130_fd_sc_hd__nand2_2 _13063_ (.A(_03912_),
    .B(_03913_),
    .Y(_03914_));
 sky130_fd_sc_hd__a21o_4 _13064_ (.A1(_03737_),
    .A2(_03755_),
    .B1(_03914_),
    .X(_03915_));
 sky130_fd_sc_hd__nand3_2 _13065_ (.A(_03737_),
    .B(_03755_),
    .C(_03914_),
    .Y(_03916_));
 sky130_fd_sc_hd__a22oi_2 _13066_ (.A1(net328),
    .A2(net802),
    .B1(net812),
    .B2(net318),
    .Y(_03917_));
 sky130_fd_sc_hd__and4_1 _13067_ (.A(net318),
    .B(net328),
    .C(net802),
    .D(net812),
    .X(_03918_));
 sky130_fd_sc_hd__nor2_1 _13068_ (.A(_03917_),
    .B(_03918_),
    .Y(_03919_));
 sky130_fd_sc_hd__nand2_2 _13069_ (.A(net337),
    .B(net795),
    .Y(_03920_));
 sky130_fd_sc_hd__xnor2_2 _13070_ (.A(_03919_),
    .B(_03920_),
    .Y(_03922_));
 sky130_fd_sc_hd__o21a_2 _13071_ (.A1(_03749_),
    .A2(_03751_),
    .B1(_03922_),
    .X(_03923_));
 sky130_fd_sc_hd__nor3_1 _13072_ (.A(_03749_),
    .B(_03751_),
    .C(_03922_),
    .Y(_03924_));
 sky130_fd_sc_hd__nor2_2 _13073_ (.A(_03923_),
    .B(_03924_),
    .Y(_03925_));
 sky130_fd_sc_hd__a21o_2 _13074_ (.A1(_03915_),
    .A2(_03916_),
    .B1(_03925_),
    .X(_03926_));
 sky130_fd_sc_hd__nand3_4 _13075_ (.A(_03915_),
    .B(_03916_),
    .C(_03925_),
    .Y(_03927_));
 sky130_fd_sc_hd__o211a_2 _13076_ (.A1(_03759_),
    .A2(_03772_),
    .B1(_03926_),
    .C1(_03927_),
    .X(_03928_));
 sky130_fd_sc_hd__a211oi_4 _13077_ (.A1(_03926_),
    .A2(_03927_),
    .B1(_03759_),
    .C1(_03772_),
    .Y(_03929_));
 sky130_fd_sc_hd__a21bo_2 _13078_ (.A1(_03802_),
    .A2(_03820_),
    .B1_N(_03819_),
    .X(_03930_));
 sky130_fd_sc_hd__a22oi_4 _13079_ (.A1(net375),
    .A2(net742),
    .B1(net751),
    .B2(net366),
    .Y(_03931_));
 sky130_fd_sc_hd__and4_2 _13080_ (.A(net366),
    .B(net375),
    .C(net742),
    .D(net751),
    .X(_03933_));
 sky130_fd_sc_hd__nand2_1 _13081_ (.A(net384),
    .B(net733),
    .Y(_03934_));
 sky130_fd_sc_hd__o21a_1 _13082_ (.A1(_03931_),
    .A2(_03933_),
    .B1(_03934_),
    .X(_03935_));
 sky130_fd_sc_hd__nor3_2 _13083_ (.A(_03931_),
    .B(_03933_),
    .C(_03934_),
    .Y(_03936_));
 sky130_fd_sc_hd__nor2_2 _13084_ (.A(_03935_),
    .B(_03936_),
    .Y(_03937_));
 sky130_fd_sc_hd__or3_1 _13085_ (.A(_03782_),
    .B(_03785_),
    .C(_03937_),
    .X(_03938_));
 sky130_fd_sc_hd__o21ai_2 _13086_ (.A1(_03782_),
    .A2(_03785_),
    .B1(_03937_),
    .Y(_03939_));
 sky130_fd_sc_hd__and2_1 _13087_ (.A(_03938_),
    .B(_03939_),
    .X(_03940_));
 sky130_fd_sc_hd__nand3_2 _13088_ (.A(net393),
    .B(net725),
    .C(_03940_),
    .Y(_03941_));
 sky130_fd_sc_hd__a21o_1 _13089_ (.A1(net393),
    .A2(net725),
    .B1(_03940_),
    .X(_03942_));
 sky130_fd_sc_hd__nand2_1 _13090_ (.A(_03941_),
    .B(_03942_),
    .Y(_03944_));
 sky130_fd_sc_hd__a21oi_1 _13091_ (.A1(_03788_),
    .A2(_03791_),
    .B1(_03944_),
    .Y(_03945_));
 sky130_fd_sc_hd__and3_1 _13092_ (.A(_03788_),
    .B(_03791_),
    .C(_03944_),
    .X(_03946_));
 sky130_fd_sc_hd__nor2_1 _13093_ (.A(_03945_),
    .B(_03946_),
    .Y(_03947_));
 sky130_fd_sc_hd__nand2_1 _13094_ (.A(net401),
    .B(net715),
    .Y(_03948_));
 sky130_fd_sc_hd__xnor2_1 _13095_ (.A(_03947_),
    .B(_03948_),
    .Y(_03949_));
 sky130_fd_sc_hd__o21ba_1 _13096_ (.A1(_03760_),
    .A2(_03763_),
    .B1_N(_03761_),
    .X(_03950_));
 sky130_fd_sc_hd__a22oi_2 _13097_ (.A1(net352),
    .A2(net773),
    .B1(net779),
    .B2(net344),
    .Y(_03951_));
 sky130_fd_sc_hd__and4_1 _13098_ (.A(net344),
    .B(net352),
    .C(net773),
    .D(net779),
    .X(_03952_));
 sky130_fd_sc_hd__nor2_1 _13099_ (.A(_03951_),
    .B(_03952_),
    .Y(_03953_));
 sky130_fd_sc_hd__nand2_2 _13100_ (.A(net359),
    .B(net761),
    .Y(_03955_));
 sky130_fd_sc_hd__xnor2_2 _13101_ (.A(_03953_),
    .B(_03955_),
    .Y(_03956_));
 sky130_fd_sc_hd__and2b_1 _13102_ (.A_N(_03950_),
    .B(_03956_),
    .X(_03957_));
 sky130_fd_sc_hd__xnor2_1 _13103_ (.A(_03950_),
    .B(_03956_),
    .Y(_03958_));
 sky130_fd_sc_hd__o21ba_1 _13104_ (.A1(_03804_),
    .A2(_03807_),
    .B1_N(_03805_),
    .X(_03959_));
 sky130_fd_sc_hd__and2b_1 _13105_ (.A_N(_03959_),
    .B(_03958_),
    .X(_03960_));
 sky130_fd_sc_hd__xor2_1 _13106_ (.A(_03958_),
    .B(_03959_),
    .X(_03961_));
 sky130_fd_sc_hd__nor2_1 _13107_ (.A(_03809_),
    .B(_03813_),
    .Y(_03962_));
 sky130_fd_sc_hd__or2_4 _13108_ (.A(_03961_),
    .B(_03962_),
    .X(_03963_));
 sky130_fd_sc_hd__nand2_1 _13109_ (.A(_03961_),
    .B(_03962_),
    .Y(_03964_));
 sky130_fd_sc_hd__and2_1 _13110_ (.A(_03963_),
    .B(_03964_),
    .X(_03966_));
 sky130_fd_sc_hd__and2b_2 _13111_ (.A_N(_03816_),
    .B(_03966_),
    .X(_03967_));
 sky130_fd_sc_hd__xnor2_1 _13112_ (.A(_03816_),
    .B(_03966_),
    .Y(_03968_));
 sky130_fd_sc_hd__and2_2 _13113_ (.A(_03949_),
    .B(_03968_),
    .X(_03969_));
 sky130_fd_sc_hd__nor2_1 _13114_ (.A(_03949_),
    .B(_03968_),
    .Y(_03970_));
 sky130_fd_sc_hd__or2_1 _13115_ (.A(_03969_),
    .B(_03970_),
    .X(_03971_));
 sky130_fd_sc_hd__a21o_1 _13116_ (.A1(_03765_),
    .A2(_03769_),
    .B1(_03971_),
    .X(_03972_));
 sky130_fd_sc_hd__nand3_1 _13117_ (.A(_03765_),
    .B(_03769_),
    .C(_03971_),
    .Y(_03973_));
 sky130_fd_sc_hd__nand2_1 _13118_ (.A(_03972_),
    .B(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hd__nand2b_1 _13119_ (.A_N(_03974_),
    .B(_03930_),
    .Y(_03975_));
 sky130_fd_sc_hd__xor2_2 _13120_ (.A(_03930_),
    .B(_03974_),
    .X(_03977_));
 sky130_fd_sc_hd__nor3_2 _13121_ (.A(_03928_),
    .B(_03929_),
    .C(_03977_),
    .Y(_03978_));
 sky130_fd_sc_hd__o21a_1 _13122_ (.A1(_03928_),
    .A2(_03929_),
    .B1(_03977_),
    .X(_03979_));
 sky130_fd_sc_hd__or2_2 _13123_ (.A(_03978_),
    .B(_03979_),
    .X(_03980_));
 sky130_fd_sc_hd__a21oi_4 _13124_ (.A1(_03776_),
    .A2(_03829_),
    .B1(_03980_),
    .Y(_03981_));
 sky130_fd_sc_hd__and3_4 _13125_ (.A(_03776_),
    .B(_03829_),
    .C(_03980_),
    .X(_03982_));
 sky130_fd_sc_hd__a211oi_4 _13126_ (.A1(_03824_),
    .A2(_03826_),
    .B1(_03981_),
    .C1(_03982_),
    .Y(_03983_));
 sky130_fd_sc_hd__a211o_2 _13127_ (.A1(_03824_),
    .A2(_03826_),
    .B1(_03981_),
    .C1(_03982_),
    .X(_03984_));
 sky130_fd_sc_hd__o211ai_4 _13128_ (.A1(_03981_),
    .A2(_03982_),
    .B1(_03824_),
    .C1(_03826_),
    .Y(_03985_));
 sky130_fd_sc_hd__o211a_2 _13129_ (.A1(_03831_),
    .A2(_03833_),
    .B1(_03984_),
    .C1(_03985_),
    .X(_03986_));
 sky130_fd_sc_hd__a211oi_4 _13130_ (.A1(_03984_),
    .A2(_03985_),
    .B1(_03831_),
    .C1(_03833_),
    .Y(_03988_));
 sky130_fd_sc_hd__a211oi_4 _13131_ (.A1(_03795_),
    .A2(_03799_),
    .B1(_03986_),
    .C1(_03988_),
    .Y(_03989_));
 sky130_fd_sc_hd__o211a_1 _13132_ (.A1(_03986_),
    .A2(_03988_),
    .B1(_03795_),
    .C1(_03799_),
    .X(_03990_));
 sky130_fd_sc_hd__a211o_2 _13133_ (.A1(_03838_),
    .A2(_03842_),
    .B1(_03989_),
    .C1(_03990_),
    .X(_03991_));
 sky130_fd_sc_hd__inv_2 _13134_ (.A(_03991_),
    .Y(_03992_));
 sky130_fd_sc_hd__o211a_1 _13135_ (.A1(_03989_),
    .A2(_03990_),
    .B1(_03838_),
    .C1(_03842_),
    .X(_03993_));
 sky130_fd_sc_hd__inv_2 _13136_ (.A(_03993_),
    .Y(_03994_));
 sky130_fd_sc_hd__nand2_1 _13137_ (.A(_03991_),
    .B(_03994_),
    .Y(_03995_));
 sky130_fd_sc_hd__and2b_1 _13138_ (.A_N(_03846_),
    .B(_03857_),
    .X(_03996_));
 sky130_fd_sc_hd__or2_1 _13139_ (.A(_03995_),
    .B(_03996_),
    .X(_03997_));
 sky130_fd_sc_hd__nand2_1 _13140_ (.A(_03995_),
    .B(_03996_),
    .Y(_03999_));
 sky130_fd_sc_hd__a32o_1 _13141_ (.A1(net260),
    .A2(_03997_),
    .A3(_03999_),
    .B1(_03859_),
    .B2(_03862_),
    .X(_08682_));
 sky130_fd_sc_hd__o22a_4 _13142_ (.A1(net577),
    .A2(_02841_),
    .B1(_02856_),
    .B2(_03689_),
    .X(_04000_));
 sky130_fd_sc_hd__o21ai_2 _13143_ (.A1(net206),
    .A2(_04000_),
    .B1(net208),
    .Y(_04001_));
 sky130_fd_sc_hd__mux2_2 _13144_ (.A0(_02822_),
    .A1(_02850_),
    .S(net566),
    .X(_04002_));
 sky130_fd_sc_hd__nor2_1 _13145_ (.A(net305),
    .B(_04002_),
    .Y(_04003_));
 sky130_fd_sc_hd__a311o_1 _13146_ (.A1(net306),
    .A2(net569),
    .A3(_02830_),
    .B1(_04003_),
    .C1(net538),
    .X(_04004_));
 sky130_fd_sc_hd__a22oi_4 _13147_ (.A1(net423),
    .A2(net680),
    .B1(net698),
    .B2(net407),
    .Y(_04005_));
 sky130_fd_sc_hd__and4_1 _13148_ (.A(net407),
    .B(net423),
    .C(net680),
    .D(net698),
    .X(_04006_));
 sky130_fd_sc_hd__nor2_2 _13149_ (.A(_04005_),
    .B(_04006_),
    .Y(_04007_));
 sky130_fd_sc_hd__nand2_4 _13150_ (.A(net416),
    .B(net690),
    .Y(_04009_));
 sky130_fd_sc_hd__xnor2_4 _13151_ (.A(_04007_),
    .B(_04009_),
    .Y(_04010_));
 sky130_fd_sc_hd__o21ba_2 _13152_ (.A1(_03863_),
    .A2(_03867_),
    .B1_N(_03864_),
    .X(_04011_));
 sky130_fd_sc_hd__nand2b_2 _13153_ (.A_N(_04011_),
    .B(_04010_),
    .Y(_04012_));
 sky130_fd_sc_hd__xnor2_4 _13154_ (.A(_04010_),
    .B(_04011_),
    .Y(_04013_));
 sky130_fd_sc_hd__a22oi_2 _13155_ (.A1(net442),
    .A2(net662),
    .B1(net671),
    .B2(net432),
    .Y(_04014_));
 sky130_fd_sc_hd__and4_1 _13156_ (.A(net432),
    .B(net442),
    .C(net662),
    .D(net671),
    .X(_04015_));
 sky130_fd_sc_hd__nor2_2 _13157_ (.A(_04014_),
    .B(_04015_),
    .Y(_04016_));
 sky130_fd_sc_hd__nand2_1 _13158_ (.A(net450),
    .B(net654),
    .Y(_04017_));
 sky130_fd_sc_hd__xnor2_2 _13159_ (.A(_04016_),
    .B(_04017_),
    .Y(_04018_));
 sky130_fd_sc_hd__nand2_4 _13160_ (.A(_04013_),
    .B(_04018_),
    .Y(_04020_));
 sky130_fd_sc_hd__or2_1 _13161_ (.A(_04013_),
    .B(_04018_),
    .X(_04021_));
 sky130_fd_sc_hd__nand2_2 _13162_ (.A(_04020_),
    .B(_04021_),
    .Y(_04022_));
 sky130_fd_sc_hd__a21o_2 _13163_ (.A1(_03870_),
    .A2(_03878_),
    .B1(_04022_),
    .X(_04023_));
 sky130_fd_sc_hd__inv_2 _13164_ (.A(_04023_),
    .Y(_04024_));
 sky130_fd_sc_hd__nand3_4 _13165_ (.A(_03870_),
    .B(_03878_),
    .C(_04022_),
    .Y(_04025_));
 sky130_fd_sc_hd__o21ba_4 _13166_ (.A1(_03882_),
    .A2(_03885_),
    .B1_N(_03883_),
    .X(_04026_));
 sky130_fd_sc_hd__o21ba_4 _13167_ (.A1(_03872_),
    .A2(_03875_),
    .B1_N(_03873_),
    .X(_04027_));
 sky130_fd_sc_hd__a22oi_4 _13168_ (.A1(net470),
    .A2(net636),
    .B1(net644),
    .B2(net459),
    .Y(_04028_));
 sky130_fd_sc_hd__and4_1 _13169_ (.A(net460),
    .B(net469),
    .C(net636),
    .D(net644),
    .X(_04029_));
 sky130_fd_sc_hd__nor2_2 _13170_ (.A(_04028_),
    .B(_04029_),
    .Y(_04031_));
 sky130_fd_sc_hd__nand2_4 _13171_ (.A(net479),
    .B(net627),
    .Y(_04032_));
 sky130_fd_sc_hd__xnor2_4 _13172_ (.A(_04031_),
    .B(_04032_),
    .Y(_04033_));
 sky130_fd_sc_hd__and2b_2 _13173_ (.A_N(_04027_),
    .B(_04033_),
    .X(_04034_));
 sky130_fd_sc_hd__xnor2_4 _13174_ (.A(_04027_),
    .B(_04033_),
    .Y(_04035_));
 sky130_fd_sc_hd__and2b_1 _13175_ (.A_N(_04026_),
    .B(_04035_),
    .X(_04036_));
 sky130_fd_sc_hd__xnor2_4 _13176_ (.A(_04026_),
    .B(_04035_),
    .Y(_04037_));
 sky130_fd_sc_hd__a21oi_4 _13177_ (.A1(_04023_),
    .A2(_04025_),
    .B1(_04037_),
    .Y(_04038_));
 sky130_fd_sc_hd__and3_4 _13178_ (.A(_04023_),
    .B(_04025_),
    .C(_04037_),
    .X(_04039_));
 sky130_fd_sc_hd__a211o_4 _13179_ (.A1(_03880_),
    .A2(_03895_),
    .B1(_04038_),
    .C1(_04039_),
    .X(_04040_));
 sky130_fd_sc_hd__o211ai_4 _13180_ (.A1(_04038_),
    .A2(_04039_),
    .B1(_03880_),
    .C1(_03895_),
    .Y(_04042_));
 sky130_fd_sc_hd__nand2_1 _13181_ (.A(_03887_),
    .B(_03891_),
    .Y(_04043_));
 sky130_fd_sc_hd__and3_1 _13182_ (.A(net485),
    .B(net619),
    .C(_03740_),
    .X(_04044_));
 sky130_fd_sc_hd__and2_1 _13183_ (.A(_04043_),
    .B(_04044_),
    .X(_04045_));
 sky130_fd_sc_hd__xnor2_1 _13184_ (.A(_04043_),
    .B(_04044_),
    .Y(_04046_));
 sky130_fd_sc_hd__nor2_2 _13185_ (.A(_03904_),
    .B(_04046_),
    .Y(_04047_));
 sky130_fd_sc_hd__and2_1 _13186_ (.A(_03904_),
    .B(_04046_),
    .X(_04048_));
 sky130_fd_sc_hd__nor2_4 _13187_ (.A(_04047_),
    .B(_04048_),
    .Y(_04049_));
 sky130_fd_sc_hd__and3_2 _13188_ (.A(_04040_),
    .B(_04042_),
    .C(_04049_),
    .X(_04050_));
 sky130_fd_sc_hd__nand3_4 _13189_ (.A(_04040_),
    .B(_04042_),
    .C(_04049_),
    .Y(_04051_));
 sky130_fd_sc_hd__a21oi_4 _13190_ (.A1(_04040_),
    .A2(_04042_),
    .B1(_04049_),
    .Y(_04053_));
 sky130_fd_sc_hd__a211o_4 _13191_ (.A1(_03897_),
    .A2(_03912_),
    .B1(_04050_),
    .C1(_04053_),
    .X(_04054_));
 sky130_fd_sc_hd__o211ai_4 _13192_ (.A1(_04050_),
    .A2(_04053_),
    .B1(_03897_),
    .C1(_03912_),
    .Y(_04055_));
 sky130_fd_sc_hd__a22oi_4 _13193_ (.A1(net328),
    .A2(net799),
    .B1(net802),
    .B2(net318),
    .Y(_04056_));
 sky130_fd_sc_hd__and4_1 _13194_ (.A(net324),
    .B(net334),
    .C(net795),
    .D(net802),
    .X(_04057_));
 sky130_fd_sc_hd__nor2_1 _13195_ (.A(_04056_),
    .B(_04057_),
    .Y(_04058_));
 sky130_fd_sc_hd__nand2_2 _13196_ (.A(net337),
    .B(net779),
    .Y(_04059_));
 sky130_fd_sc_hd__xnor2_2 _13197_ (.A(_04058_),
    .B(_04059_),
    .Y(_04060_));
 sky130_fd_sc_hd__o21a_2 _13198_ (.A1(_03906_),
    .A2(_03909_),
    .B1(_04060_),
    .X(_04061_));
 sky130_fd_sc_hd__nor3_1 _13199_ (.A(_03906_),
    .B(_03909_),
    .C(_04060_),
    .Y(_04062_));
 sky130_fd_sc_hd__nor2_2 _13200_ (.A(_04061_),
    .B(_04062_),
    .Y(_04064_));
 sky130_fd_sc_hd__a21oi_4 _13201_ (.A1(_04054_),
    .A2(_04055_),
    .B1(_04064_),
    .Y(_04065_));
 sky130_fd_sc_hd__and3_4 _13202_ (.A(_04054_),
    .B(_04055_),
    .C(_04064_),
    .X(_04066_));
 sky130_fd_sc_hd__inv_2 _13203_ (.A(_04066_),
    .Y(_04067_));
 sky130_fd_sc_hd__a211o_4 _13204_ (.A1(_03915_),
    .A2(_03927_),
    .B1(_04065_),
    .C1(_04066_),
    .X(_04068_));
 sky130_fd_sc_hd__o211ai_4 _13205_ (.A1(_04065_),
    .A2(_04066_),
    .B1(_03915_),
    .C1(_03927_),
    .Y(_04069_));
 sky130_fd_sc_hd__nand2_4 _13206_ (.A(net401),
    .B(net708),
    .Y(_04070_));
 sky130_fd_sc_hd__a22oi_4 _13207_ (.A1(net375),
    .A2(net733),
    .B1(net742),
    .B2(net366),
    .Y(_04071_));
 sky130_fd_sc_hd__and4_2 _13208_ (.A(net366),
    .B(net375),
    .C(net733),
    .D(net742),
    .X(_04072_));
 sky130_fd_sc_hd__nand2_1 _13209_ (.A(net384),
    .B(net725),
    .Y(_04073_));
 sky130_fd_sc_hd__o21a_1 _13210_ (.A1(_04071_),
    .A2(_04072_),
    .B1(_04073_),
    .X(_04075_));
 sky130_fd_sc_hd__nor3_2 _13211_ (.A(_04071_),
    .B(_04072_),
    .C(_04073_),
    .Y(_04076_));
 sky130_fd_sc_hd__nor2_1 _13212_ (.A(_04075_),
    .B(_04076_),
    .Y(_04077_));
 sky130_fd_sc_hd__or3_1 _13213_ (.A(_03933_),
    .B(_03936_),
    .C(_04077_),
    .X(_04078_));
 sky130_fd_sc_hd__o21ai_1 _13214_ (.A1(_03933_),
    .A2(_03936_),
    .B1(_04077_),
    .Y(_04079_));
 sky130_fd_sc_hd__and2_1 _13215_ (.A(_04078_),
    .B(_04079_),
    .X(_04080_));
 sky130_fd_sc_hd__nand3_1 _13216_ (.A(net392),
    .B(net715),
    .C(_04080_),
    .Y(_04081_));
 sky130_fd_sc_hd__a21o_1 _13217_ (.A1(net392),
    .A2(net715),
    .B1(_04080_),
    .X(_04082_));
 sky130_fd_sc_hd__nand2_1 _13218_ (.A(_04081_),
    .B(_04082_),
    .Y(_04083_));
 sky130_fd_sc_hd__a21o_2 _13219_ (.A1(_03939_),
    .A2(_03941_),
    .B1(_04083_),
    .X(_04084_));
 sky130_fd_sc_hd__nand3_1 _13220_ (.A(_03939_),
    .B(_03941_),
    .C(_04083_),
    .Y(_04086_));
 sky130_fd_sc_hd__nand2_1 _13221_ (.A(_04084_),
    .B(_04086_),
    .Y(_04087_));
 sky130_fd_sc_hd__or2_2 _13222_ (.A(_04070_),
    .B(_04087_),
    .X(_04088_));
 sky130_fd_sc_hd__nand2_1 _13223_ (.A(_04070_),
    .B(_04087_),
    .Y(_04089_));
 sky130_fd_sc_hd__and2_2 _13224_ (.A(_04088_),
    .B(_04089_),
    .X(_04090_));
 sky130_fd_sc_hd__o21ba_1 _13225_ (.A1(_03917_),
    .A2(_03920_),
    .B1_N(_03918_),
    .X(_04091_));
 sky130_fd_sc_hd__a22oi_2 _13226_ (.A1(net352),
    .A2(net761),
    .B1(net773),
    .B2(net344),
    .Y(_04092_));
 sky130_fd_sc_hd__and4_1 _13227_ (.A(net344),
    .B(net352),
    .C(net761),
    .D(net773),
    .X(_04093_));
 sky130_fd_sc_hd__nor2_1 _13228_ (.A(_04092_),
    .B(_04093_),
    .Y(_04094_));
 sky130_fd_sc_hd__nand2_2 _13229_ (.A(net359),
    .B(net751),
    .Y(_04095_));
 sky130_fd_sc_hd__xnor2_2 _13230_ (.A(_04094_),
    .B(_04095_),
    .Y(_04097_));
 sky130_fd_sc_hd__and2b_1 _13231_ (.A_N(_04091_),
    .B(_04097_),
    .X(_04098_));
 sky130_fd_sc_hd__xnor2_1 _13232_ (.A(_04091_),
    .B(_04097_),
    .Y(_04099_));
 sky130_fd_sc_hd__o21ba_1 _13233_ (.A1(_03951_),
    .A2(_03955_),
    .B1_N(_03952_),
    .X(_04100_));
 sky130_fd_sc_hd__and2b_1 _13234_ (.A_N(_04100_),
    .B(_04099_),
    .X(_04101_));
 sky130_fd_sc_hd__xor2_1 _13235_ (.A(_04099_),
    .B(_04100_),
    .X(_04102_));
 sky130_fd_sc_hd__nor2_1 _13236_ (.A(_03957_),
    .B(_03960_),
    .Y(_04103_));
 sky130_fd_sc_hd__or2_2 _13237_ (.A(_04102_),
    .B(_04103_),
    .X(_04104_));
 sky130_fd_sc_hd__nand2_1 _13238_ (.A(_04102_),
    .B(_04103_),
    .Y(_04105_));
 sky130_fd_sc_hd__and2_2 _13239_ (.A(_04104_),
    .B(_04105_),
    .X(_04106_));
 sky130_fd_sc_hd__nand2b_2 _13240_ (.A_N(_03963_),
    .B(_04106_),
    .Y(_04108_));
 sky130_fd_sc_hd__xnor2_4 _13241_ (.A(_03963_),
    .B(_04106_),
    .Y(_04109_));
 sky130_fd_sc_hd__nand2_4 _13242_ (.A(_04090_),
    .B(_04109_),
    .Y(_04110_));
 sky130_fd_sc_hd__or2_2 _13243_ (.A(_04090_),
    .B(_04109_),
    .X(_04111_));
 sky130_fd_sc_hd__nand3_4 _13244_ (.A(_03923_),
    .B(_04110_),
    .C(_04111_),
    .Y(_04112_));
 sky130_fd_sc_hd__a21o_1 _13245_ (.A1(_04110_),
    .A2(_04111_),
    .B1(_03923_),
    .X(_04113_));
 sky130_fd_sc_hd__and2_1 _13246_ (.A(_04112_),
    .B(_04113_),
    .X(_04114_));
 sky130_fd_sc_hd__o21ai_4 _13247_ (.A1(_03967_),
    .A2(_03969_),
    .B1(_04114_),
    .Y(_04115_));
 sky130_fd_sc_hd__or3_2 _13248_ (.A(_03967_),
    .B(_03969_),
    .C(_04114_),
    .X(_04116_));
 sky130_fd_sc_hd__nand4_4 _13249_ (.A(_04068_),
    .B(_04069_),
    .C(_04115_),
    .D(_04116_),
    .Y(_04117_));
 sky130_fd_sc_hd__a22o_1 _13250_ (.A1(_04068_),
    .A2(_04069_),
    .B1(_04115_),
    .B2(_04116_),
    .X(_04119_));
 sky130_fd_sc_hd__o211a_1 _13251_ (.A1(_03928_),
    .A2(_03978_),
    .B1(_04117_),
    .C1(_04119_),
    .X(_04120_));
 sky130_fd_sc_hd__inv_2 _13252_ (.A(_04120_),
    .Y(_04121_));
 sky130_fd_sc_hd__a211oi_2 _13253_ (.A1(_04117_),
    .A2(_04119_),
    .B1(_03928_),
    .C1(_03978_),
    .Y(_04122_));
 sky130_fd_sc_hd__a211o_2 _13254_ (.A1(_03972_),
    .A2(_03975_),
    .B1(_04120_),
    .C1(_04122_),
    .X(_04123_));
 sky130_fd_sc_hd__o211ai_1 _13255_ (.A1(_04120_),
    .A2(_04122_),
    .B1(_03972_),
    .C1(_03975_),
    .Y(_04124_));
 sky130_fd_sc_hd__and2_2 _13256_ (.A(_04123_),
    .B(_04124_),
    .X(_04125_));
 sky130_fd_sc_hd__o21ai_4 _13257_ (.A1(_03981_),
    .A2(_03983_),
    .B1(_04125_),
    .Y(_04126_));
 sky130_fd_sc_hd__or3_2 _13258_ (.A(_03981_),
    .B(_03983_),
    .C(_04125_),
    .X(_04127_));
 sky130_fd_sc_hd__o21ba_1 _13259_ (.A1(_03946_),
    .A2(_03948_),
    .B1_N(_03945_),
    .X(_04128_));
 sky130_fd_sc_hd__inv_2 _13260_ (.A(_04128_),
    .Y(_04130_));
 sky130_fd_sc_hd__nand3_4 _13261_ (.A(_04126_),
    .B(_04127_),
    .C(_04130_),
    .Y(_04131_));
 sky130_fd_sc_hd__a21o_1 _13262_ (.A1(_04126_),
    .A2(_04127_),
    .B1(_04130_),
    .X(_04132_));
 sky130_fd_sc_hd__nand2_2 _13263_ (.A(_04131_),
    .B(_04132_),
    .Y(_04133_));
 sky130_fd_sc_hd__nor2_2 _13264_ (.A(_03986_),
    .B(_03989_),
    .Y(_04134_));
 sky130_fd_sc_hd__or2_1 _13265_ (.A(_04133_),
    .B(_04134_),
    .X(_04135_));
 sky130_fd_sc_hd__xnor2_1 _13266_ (.A(_04133_),
    .B(_04134_),
    .Y(_04136_));
 sky130_fd_sc_hd__o21a_1 _13267_ (.A1(_03846_),
    .A2(_03992_),
    .B1(_03994_),
    .X(_04137_));
 sky130_fd_sc_hd__nor2_1 _13268_ (.A(_03848_),
    .B(_03995_),
    .Y(_04138_));
 sky130_fd_sc_hd__a21oi_1 _13269_ (.A1(_03854_),
    .A2(_04138_),
    .B1(_04137_),
    .Y(_04139_));
 sky130_fd_sc_hd__nand2_1 _13270_ (.A(_04136_),
    .B(_04139_),
    .Y(_04141_));
 sky130_fd_sc_hd__or2_1 _13271_ (.A(_04136_),
    .B(_04139_),
    .X(_04142_));
 sky130_fd_sc_hd__a32o_1 _13272_ (.A1(net259),
    .A2(_04141_),
    .A3(_04142_),
    .B1(_04001_),
    .B2(_04004_),
    .X(_08683_));
 sky130_fd_sc_hd__o22a_4 _13273_ (.A1(net566),
    .A2(_03015_),
    .B1(_03021_),
    .B2(_03689_),
    .X(_04143_));
 sky130_fd_sc_hd__o21ai_1 _13274_ (.A1(net206),
    .A2(_04143_),
    .B1(net208),
    .Y(_04144_));
 sky130_fd_sc_hd__mux2_2 _13275_ (.A0(_03006_),
    .A1(_03018_),
    .S(net567),
    .X(_04145_));
 sky130_fd_sc_hd__nor2_1 _13276_ (.A(net305),
    .B(_04145_),
    .Y(_04146_));
 sky130_fd_sc_hd__a311o_1 _13277_ (.A1(net306),
    .A2(net570),
    .A3(_03010_),
    .B1(_04146_),
    .C1(net539),
    .X(_04147_));
 sky130_fd_sc_hd__a22oi_4 _13278_ (.A1(net423),
    .A2(net670),
    .B1(net689),
    .B2(net407),
    .Y(_04148_));
 sky130_fd_sc_hd__and4_2 _13279_ (.A(net410),
    .B(net425),
    .C(net670),
    .D(net689),
    .X(_04149_));
 sky130_fd_sc_hd__nor2_4 _13280_ (.A(_04148_),
    .B(_04149_),
    .Y(_04151_));
 sky130_fd_sc_hd__nand2_2 _13281_ (.A(net416),
    .B(net680),
    .Y(_04152_));
 sky130_fd_sc_hd__xnor2_4 _13282_ (.A(_04151_),
    .B(_04152_),
    .Y(_04153_));
 sky130_fd_sc_hd__o21ba_1 _13283_ (.A1(_04005_),
    .A2(_04009_),
    .B1_N(_04006_),
    .X(_04154_));
 sky130_fd_sc_hd__nand2b_2 _13284_ (.A_N(_04154_),
    .B(_04153_),
    .Y(_04155_));
 sky130_fd_sc_hd__xnor2_1 _13285_ (.A(_04153_),
    .B(_04154_),
    .Y(_04156_));
 sky130_fd_sc_hd__a22oi_2 _13286_ (.A1(net443),
    .A2(net654),
    .B1(net662),
    .B2(net432),
    .Y(_04157_));
 sky130_fd_sc_hd__and4_2 _13287_ (.A(net433),
    .B(net443),
    .C(net654),
    .D(net662),
    .X(_04158_));
 sky130_fd_sc_hd__and4bb_2 _13288_ (.A_N(_04157_),
    .B_N(_04158_),
    .C(net450),
    .D(net644),
    .X(_04159_));
 sky130_fd_sc_hd__o2bb2a_1 _13289_ (.A1_N(net450),
    .A2_N(net644),
    .B1(_04157_),
    .B2(_04158_),
    .X(_04160_));
 sky130_fd_sc_hd__nor2_1 _13290_ (.A(_04159_),
    .B(_04160_),
    .Y(_04162_));
 sky130_fd_sc_hd__nand2_2 _13291_ (.A(_04156_),
    .B(_04162_),
    .Y(_04163_));
 sky130_fd_sc_hd__or2_1 _13292_ (.A(_04156_),
    .B(_04162_),
    .X(_04164_));
 sky130_fd_sc_hd__nand2_2 _13293_ (.A(_04163_),
    .B(_04164_),
    .Y(_04165_));
 sky130_fd_sc_hd__a21o_4 _13294_ (.A1(_04012_),
    .A2(_04020_),
    .B1(_04165_),
    .X(_04166_));
 sky130_fd_sc_hd__nand3_4 _13295_ (.A(_04012_),
    .B(_04020_),
    .C(_04165_),
    .Y(_04167_));
 sky130_fd_sc_hd__o21ba_4 _13296_ (.A1(_04028_),
    .A2(_04032_),
    .B1_N(_04029_),
    .X(_04168_));
 sky130_fd_sc_hd__a31o_4 _13297_ (.A1(net450),
    .A2(net654),
    .A3(_04016_),
    .B1(_04015_),
    .X(_04169_));
 sky130_fd_sc_hd__nand2_1 _13298_ (.A(net469),
    .B(net632),
    .Y(_04170_));
 sky130_fd_sc_hd__a21boi_2 _13299_ (.A1(net459),
    .A2(net635),
    .B1_N(_04170_),
    .Y(_04171_));
 sky130_fd_sc_hd__and4_1 _13300_ (.A(net459),
    .B(net469),
    .C(net627),
    .D(net636),
    .X(_04173_));
 sky130_fd_sc_hd__nor2_2 _13301_ (.A(_04171_),
    .B(_04173_),
    .Y(_04174_));
 sky130_fd_sc_hd__nand2_4 _13302_ (.A(net479),
    .B(net619),
    .Y(_04175_));
 sky130_fd_sc_hd__xnor2_4 _13303_ (.A(_04174_),
    .B(_04175_),
    .Y(_04176_));
 sky130_fd_sc_hd__xor2_4 _13304_ (.A(_04169_),
    .B(_04176_),
    .X(_04177_));
 sky130_fd_sc_hd__nand2b_1 _13305_ (.A_N(_04168_),
    .B(_04177_),
    .Y(_04178_));
 sky130_fd_sc_hd__xnor2_4 _13306_ (.A(_04168_),
    .B(_04177_),
    .Y(_04179_));
 sky130_fd_sc_hd__a21o_1 _13307_ (.A1(_04166_),
    .A2(_04167_),
    .B1(_04179_),
    .X(_04180_));
 sky130_fd_sc_hd__nand3_4 _13308_ (.A(_04166_),
    .B(_04167_),
    .C(_04179_),
    .Y(_04181_));
 sky130_fd_sc_hd__and2_2 _13309_ (.A(_04180_),
    .B(_04181_),
    .X(_04182_));
 sky130_fd_sc_hd__o21ai_4 _13310_ (.A1(_04024_),
    .A2(_04039_),
    .B1(_04182_),
    .Y(_04184_));
 sky130_fd_sc_hd__inv_2 _13311_ (.A(_04184_),
    .Y(_04185_));
 sky130_fd_sc_hd__or3_4 _13312_ (.A(_04024_),
    .B(_04039_),
    .C(_04182_),
    .X(_04186_));
 sky130_fd_sc_hd__o21ai_4 _13313_ (.A1(_04034_),
    .A2(_04036_),
    .B1(_03901_),
    .Y(_04187_));
 sky130_fd_sc_hd__or3_1 _13314_ (.A(_03901_),
    .B(_04034_),
    .C(_04036_),
    .X(_04188_));
 sky130_fd_sc_hd__and2_2 _13315_ (.A(_04187_),
    .B(_04188_),
    .X(_04189_));
 sky130_fd_sc_hd__a21oi_4 _13316_ (.A1(_04184_),
    .A2(_04186_),
    .B1(_04189_),
    .Y(_04190_));
 sky130_fd_sc_hd__and3_4 _13317_ (.A(_04184_),
    .B(_04186_),
    .C(_04189_),
    .X(_04191_));
 sky130_fd_sc_hd__a211o_4 _13318_ (.A1(_04040_),
    .A2(_04051_),
    .B1(_04190_),
    .C1(_04191_),
    .X(_04192_));
 sky130_fd_sc_hd__o211ai_4 _13319_ (.A1(_04190_),
    .A2(_04191_),
    .B1(_04040_),
    .C1(_04051_),
    .Y(_04193_));
 sky130_fd_sc_hd__a22oi_2 _13320_ (.A1(net333),
    .A2(net787),
    .B1(net795),
    .B2(net323),
    .Y(_04195_));
 sky130_fd_sc_hd__and4_1 _13321_ (.A(net323),
    .B(net333),
    .C(net779),
    .D(net795),
    .X(_04196_));
 sky130_fd_sc_hd__nor2_1 _13322_ (.A(_04195_),
    .B(_04196_),
    .Y(_04197_));
 sky130_fd_sc_hd__nand2_2 _13323_ (.A(net338),
    .B(net776),
    .Y(_04198_));
 sky130_fd_sc_hd__xnor2_2 _13324_ (.A(_04197_),
    .B(_04198_),
    .Y(_04199_));
 sky130_fd_sc_hd__o21a_2 _13325_ (.A1(_04045_),
    .A2(_04047_),
    .B1(_04199_),
    .X(_04200_));
 sky130_fd_sc_hd__nor3_1 _13326_ (.A(_04045_),
    .B(_04047_),
    .C(_04199_),
    .Y(_04201_));
 sky130_fd_sc_hd__nor2_2 _13327_ (.A(_04200_),
    .B(_04201_),
    .Y(_04202_));
 sky130_fd_sc_hd__a21o_1 _13328_ (.A1(_04192_),
    .A2(_04193_),
    .B1(_04202_),
    .X(_04203_));
 sky130_fd_sc_hd__nand3_4 _13329_ (.A(_04192_),
    .B(_04193_),
    .C(_04202_),
    .Y(_04204_));
 sky130_fd_sc_hd__nand2_2 _13330_ (.A(_04203_),
    .B(_04204_),
    .Y(_04206_));
 sky130_fd_sc_hd__a21oi_4 _13331_ (.A1(_04054_),
    .A2(_04067_),
    .B1(_04206_),
    .Y(_04207_));
 sky130_fd_sc_hd__and3_2 _13332_ (.A(_04054_),
    .B(_04067_),
    .C(_04206_),
    .X(_04208_));
 sky130_fd_sc_hd__a22oi_4 _13333_ (.A1(net375),
    .A2(net725),
    .B1(net733),
    .B2(net366),
    .Y(_04209_));
 sky130_fd_sc_hd__and4_2 _13334_ (.A(net366),
    .B(net375),
    .C(net725),
    .D(net733),
    .X(_04210_));
 sky130_fd_sc_hd__nand2_1 _13335_ (.A(net384),
    .B(net715),
    .Y(_04211_));
 sky130_fd_sc_hd__o21a_1 _13336_ (.A1(_04209_),
    .A2(_04210_),
    .B1(_04211_),
    .X(_04212_));
 sky130_fd_sc_hd__nor3_2 _13337_ (.A(_04209_),
    .B(_04210_),
    .C(_04211_),
    .Y(_04213_));
 sky130_fd_sc_hd__nor2_1 _13338_ (.A(_04212_),
    .B(_04213_),
    .Y(_04214_));
 sky130_fd_sc_hd__or3_1 _13339_ (.A(_04072_),
    .B(_04076_),
    .C(_04214_),
    .X(_04215_));
 sky130_fd_sc_hd__o21ai_2 _13340_ (.A1(_04072_),
    .A2(_04076_),
    .B1(_04214_),
    .Y(_04217_));
 sky130_fd_sc_hd__and2_1 _13341_ (.A(_04215_),
    .B(_04217_),
    .X(_04218_));
 sky130_fd_sc_hd__nand3_2 _13342_ (.A(net392),
    .B(net706),
    .C(_04218_),
    .Y(_04219_));
 sky130_fd_sc_hd__a21o_1 _13343_ (.A1(net392),
    .A2(net706),
    .B1(_04218_),
    .X(_04220_));
 sky130_fd_sc_hd__nand2_1 _13344_ (.A(_04219_),
    .B(_04220_),
    .Y(_04221_));
 sky130_fd_sc_hd__a21oi_1 _13345_ (.A1(_04079_),
    .A2(_04081_),
    .B1(_04221_),
    .Y(_04222_));
 sky130_fd_sc_hd__and3_1 _13346_ (.A(_04079_),
    .B(_04081_),
    .C(_04221_),
    .X(_04223_));
 sky130_fd_sc_hd__nor2_1 _13347_ (.A(_04222_),
    .B(_04223_),
    .Y(_04224_));
 sky130_fd_sc_hd__nand2_2 _13348_ (.A(net400),
    .B(net699),
    .Y(_04225_));
 sky130_fd_sc_hd__xnor2_2 _13349_ (.A(_04224_),
    .B(_04225_),
    .Y(_04226_));
 sky130_fd_sc_hd__o21ba_4 _13350_ (.A1(_04056_),
    .A2(_04059_),
    .B1_N(_04057_),
    .X(_04228_));
 sky130_fd_sc_hd__a22oi_4 _13351_ (.A1(net351),
    .A2(net752),
    .B1(net765),
    .B2(net345),
    .Y(_04229_));
 sky130_fd_sc_hd__and4_1 _13352_ (.A(net345),
    .B(net351),
    .C(net752),
    .D(net761),
    .X(_04230_));
 sky130_fd_sc_hd__nor2_2 _13353_ (.A(_04229_),
    .B(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__nand2_4 _13354_ (.A(net359),
    .B(net742),
    .Y(_04232_));
 sky130_fd_sc_hd__xnor2_4 _13355_ (.A(_04231_),
    .B(_04232_),
    .Y(_04233_));
 sky130_fd_sc_hd__and2b_1 _13356_ (.A_N(_04228_),
    .B(_04233_),
    .X(_04234_));
 sky130_fd_sc_hd__xnor2_4 _13357_ (.A(_04228_),
    .B(_04233_),
    .Y(_04235_));
 sky130_fd_sc_hd__o21ba_2 _13358_ (.A1(_04092_),
    .A2(_04095_),
    .B1_N(_04093_),
    .X(_04236_));
 sky130_fd_sc_hd__and2b_1 _13359_ (.A_N(_04236_),
    .B(_04235_),
    .X(_04237_));
 sky130_fd_sc_hd__xor2_2 _13360_ (.A(_04235_),
    .B(_04236_),
    .X(_04239_));
 sky130_fd_sc_hd__nor2_1 _13361_ (.A(_04098_),
    .B(_04101_),
    .Y(_04240_));
 sky130_fd_sc_hd__nor2_2 _13362_ (.A(_04239_),
    .B(_04240_),
    .Y(_04241_));
 sky130_fd_sc_hd__and2_1 _13363_ (.A(_04239_),
    .B(_04240_),
    .X(_04242_));
 sky130_fd_sc_hd__nor2_2 _13364_ (.A(_04241_),
    .B(_04242_),
    .Y(_04243_));
 sky130_fd_sc_hd__nand2b_2 _13365_ (.A_N(_04104_),
    .B(_04243_),
    .Y(_04244_));
 sky130_fd_sc_hd__xnor2_2 _13366_ (.A(_04104_),
    .B(_04243_),
    .Y(_04245_));
 sky130_fd_sc_hd__nand2_4 _13367_ (.A(_04226_),
    .B(_04245_),
    .Y(_04246_));
 sky130_fd_sc_hd__or2_2 _13368_ (.A(_04226_),
    .B(_04245_),
    .X(_04247_));
 sky130_fd_sc_hd__and3_2 _13369_ (.A(_04061_),
    .B(_04246_),
    .C(_04247_),
    .X(_04248_));
 sky130_fd_sc_hd__a21oi_4 _13370_ (.A1(_04246_),
    .A2(_04247_),
    .B1(_04061_),
    .Y(_04250_));
 sky130_fd_sc_hd__a211oi_4 _13371_ (.A1(_04108_),
    .A2(_04110_),
    .B1(_04248_),
    .C1(_04250_),
    .Y(_04251_));
 sky130_fd_sc_hd__o211a_2 _13372_ (.A1(_04248_),
    .A2(_04250_),
    .B1(_04108_),
    .C1(_04110_),
    .X(_04252_));
 sky130_fd_sc_hd__nor4_4 _13373_ (.A(_04207_),
    .B(_04208_),
    .C(_04251_),
    .D(_04252_),
    .Y(_04253_));
 sky130_fd_sc_hd__o22a_2 _13374_ (.A1(_04207_),
    .A2(_04208_),
    .B1(_04251_),
    .B2(_04252_),
    .X(_04254_));
 sky130_fd_sc_hd__a211oi_4 _13375_ (.A1(_04068_),
    .A2(_04117_),
    .B1(_04253_),
    .C1(_04254_),
    .Y(_04255_));
 sky130_fd_sc_hd__o211a_2 _13376_ (.A1(_04253_),
    .A2(_04254_),
    .B1(_04068_),
    .C1(_04117_),
    .X(_04256_));
 sky130_fd_sc_hd__a211oi_4 _13377_ (.A1(_04112_),
    .A2(_04115_),
    .B1(_04255_),
    .C1(_04256_),
    .Y(_04257_));
 sky130_fd_sc_hd__o211a_2 _13378_ (.A1(_04255_),
    .A2(_04256_),
    .B1(_04112_),
    .C1(_04115_),
    .X(_04258_));
 sky130_fd_sc_hd__a211oi_4 _13379_ (.A1(_04121_),
    .A2(_04123_),
    .B1(_04257_),
    .C1(_04258_),
    .Y(_04259_));
 sky130_fd_sc_hd__o211a_2 _13380_ (.A1(_04257_),
    .A2(_04258_),
    .B1(_04121_),
    .C1(_04123_),
    .X(_04261_));
 sky130_fd_sc_hd__a211oi_4 _13381_ (.A1(_04084_),
    .A2(_04088_),
    .B1(_04259_),
    .C1(_04261_),
    .Y(_04262_));
 sky130_fd_sc_hd__o211a_2 _13382_ (.A1(_04259_),
    .A2(_04261_),
    .B1(_04084_),
    .C1(_04088_),
    .X(_04263_));
 sky130_fd_sc_hd__o211a_2 _13383_ (.A1(_04262_),
    .A2(_04263_),
    .B1(_04126_),
    .C1(_04131_),
    .X(_04264_));
 sky130_fd_sc_hd__a211oi_4 _13384_ (.A1(_04126_),
    .A2(_04131_),
    .B1(_04262_),
    .C1(_04263_),
    .Y(_04265_));
 sky130_fd_sc_hd__nor2_1 _13385_ (.A(_04264_),
    .B(_04265_),
    .Y(_04266_));
 sky130_fd_sc_hd__nand2_1 _13386_ (.A(_04135_),
    .B(_04142_),
    .Y(_04267_));
 sky130_fd_sc_hd__nand2_1 _13387_ (.A(_04266_),
    .B(_04267_),
    .Y(_04268_));
 sky130_fd_sc_hd__or2_1 _13388_ (.A(_04266_),
    .B(_04267_),
    .X(_04269_));
 sky130_fd_sc_hd__a32o_1 _13389_ (.A1(net259),
    .A2(_04268_),
    .A3(_04269_),
    .B1(_04144_),
    .B2(_04147_),
    .X(_08654_));
 sky130_fd_sc_hd__mux2_4 _13390_ (.A0(_03176_),
    .A1(_03192_),
    .S(net568),
    .X(_04271_));
 sky130_fd_sc_hd__o21ai_2 _13391_ (.A1(net206),
    .A2(_04271_),
    .B1(net208),
    .Y(_04272_));
 sky130_fd_sc_hd__mux2_1 _13392_ (.A0(_03179_),
    .A1(_03184_),
    .S(net300),
    .X(_04273_));
 sky130_fd_sc_hd__nor2_1 _13393_ (.A(net305),
    .B(_04273_),
    .Y(_04274_));
 sky130_fd_sc_hd__a311o_1 _13394_ (.A1(net305),
    .A2(net569),
    .A3(_03186_),
    .B1(_04274_),
    .C1(net538),
    .X(_04275_));
 sky130_fd_sc_hd__a22o_2 _13395_ (.A1(net425),
    .A2(net663),
    .B1(net680),
    .B2(net407),
    .X(_04276_));
 sky130_fd_sc_hd__nand4_4 _13396_ (.A(net407),
    .B(net425),
    .C(net663),
    .D(net680),
    .Y(_04277_));
 sky130_fd_sc_hd__nand2_1 _13397_ (.A(net416),
    .B(net670),
    .Y(_04278_));
 sky130_fd_sc_hd__nand3b_4 _13398_ (.A_N(_04278_),
    .B(_04277_),
    .C(_04276_),
    .Y(_04279_));
 sky130_fd_sc_hd__a21bo_1 _13399_ (.A1(_04276_),
    .A2(_04277_),
    .B1_N(_04278_),
    .X(_04280_));
 sky130_fd_sc_hd__a31o_1 _13400_ (.A1(net416),
    .A2(net680),
    .A3(_04151_),
    .B1(_04149_),
    .X(_04282_));
 sky130_fd_sc_hd__nand3_2 _13401_ (.A(_04279_),
    .B(_04280_),
    .C(_04282_),
    .Y(_04283_));
 sky130_fd_sc_hd__a21o_2 _13402_ (.A1(_04279_),
    .A2(_04280_),
    .B1(_04282_),
    .X(_04284_));
 sky130_fd_sc_hd__nand2_2 _13403_ (.A(_04283_),
    .B(_04284_),
    .Y(_04285_));
 sky130_fd_sc_hd__a22oi_4 _13404_ (.A1(net443),
    .A2(net644),
    .B1(net654),
    .B2(net432),
    .Y(_04286_));
 sky130_fd_sc_hd__and4_2 _13405_ (.A(net433),
    .B(net443),
    .C(net644),
    .D(net654),
    .X(_04287_));
 sky130_fd_sc_hd__nor2_4 _13406_ (.A(_04286_),
    .B(_04287_),
    .Y(_04288_));
 sky130_fd_sc_hd__nand2_2 _13407_ (.A(net450),
    .B(net636),
    .Y(_04289_));
 sky130_fd_sc_hd__xnor2_4 _13408_ (.A(_04288_),
    .B(_04289_),
    .Y(_04290_));
 sky130_fd_sc_hd__xor2_4 _13409_ (.A(_04285_),
    .B(_04290_),
    .X(_04291_));
 sky130_fd_sc_hd__a21o_4 _13410_ (.A1(_04155_),
    .A2(_04163_),
    .B1(_04291_),
    .X(_04293_));
 sky130_fd_sc_hd__nand3_4 _13411_ (.A(_04155_),
    .B(_04163_),
    .C(_04291_),
    .Y(_04294_));
 sky130_fd_sc_hd__o21ba_4 _13412_ (.A1(_04171_),
    .A2(_04175_),
    .B1_N(_04173_),
    .X(_04295_));
 sky130_fd_sc_hd__a22oi_2 _13413_ (.A1(net469),
    .A2(net624),
    .B1(net627),
    .B2(net459),
    .Y(_04296_));
 sky130_fd_sc_hd__and4_1 _13414_ (.A(net459),
    .B(net469),
    .C(net624),
    .D(net632),
    .X(_04297_));
 sky130_fd_sc_hd__nor2_2 _13415_ (.A(_04296_),
    .B(_04297_),
    .Y(_04298_));
 sky130_fd_sc_hd__o21ai_4 _13416_ (.A1(_04158_),
    .A2(_04159_),
    .B1(_04298_),
    .Y(_04299_));
 sky130_fd_sc_hd__or3_1 _13417_ (.A(_04158_),
    .B(_04159_),
    .C(_04298_),
    .X(_04300_));
 sky130_fd_sc_hd__and2_2 _13418_ (.A(_04299_),
    .B(_04300_),
    .X(_04301_));
 sky130_fd_sc_hd__nand2b_2 _13419_ (.A_N(_04295_),
    .B(_04301_),
    .Y(_04302_));
 sky130_fd_sc_hd__xnor2_4 _13420_ (.A(_04295_),
    .B(_04301_),
    .Y(_04304_));
 sky130_fd_sc_hd__a21oi_4 _13421_ (.A1(_04293_),
    .A2(_04294_),
    .B1(_04304_),
    .Y(_04305_));
 sky130_fd_sc_hd__and3_2 _13422_ (.A(_04293_),
    .B(_04294_),
    .C(_04304_),
    .X(_04306_));
 sky130_fd_sc_hd__nand3_2 _13423_ (.A(_04293_),
    .B(_04294_),
    .C(_04304_),
    .Y(_04307_));
 sky130_fd_sc_hd__a211oi_4 _13424_ (.A1(_04166_),
    .A2(_04181_),
    .B1(_04305_),
    .C1(_04306_),
    .Y(_04308_));
 sky130_fd_sc_hd__clkinv_2 _13425_ (.A(_04308_),
    .Y(_04309_));
 sky130_fd_sc_hd__o211a_1 _13426_ (.A1(_04305_),
    .A2(_04306_),
    .B1(_04166_),
    .C1(_04181_),
    .X(_04310_));
 sky130_fd_sc_hd__a21bo_1 _13427_ (.A1(_04169_),
    .A2(_04176_),
    .B1_N(_04178_),
    .X(_04311_));
 sky130_fd_sc_hd__or3b_4 _13428_ (.A(_04308_),
    .B(_04310_),
    .C_N(_04311_),
    .X(_04312_));
 sky130_fd_sc_hd__o21bai_1 _13429_ (.A1(_04308_),
    .A2(_04310_),
    .B1_N(_04311_),
    .Y(_04313_));
 sky130_fd_sc_hd__and2_2 _13430_ (.A(_04312_),
    .B(_04313_),
    .X(_04315_));
 sky130_fd_sc_hd__or3_2 _13431_ (.A(_04185_),
    .B(_04191_),
    .C(_04315_),
    .X(_04316_));
 sky130_fd_sc_hd__o21ai_4 _13432_ (.A1(_04185_),
    .A2(_04191_),
    .B1(_04315_),
    .Y(_04317_));
 sky130_fd_sc_hd__a22oi_1 _13433_ (.A1(net333),
    .A2(net773),
    .B1(net779),
    .B2(net323),
    .Y(_04318_));
 sky130_fd_sc_hd__and4_1 _13434_ (.A(net323),
    .B(net333),
    .C(net773),
    .D(net779),
    .X(_04319_));
 sky130_fd_sc_hd__or2_1 _13435_ (.A(_04318_),
    .B(_04319_),
    .X(_04320_));
 sky130_fd_sc_hd__nand2_1 _13436_ (.A(net338),
    .B(net761),
    .Y(_04321_));
 sky130_fd_sc_hd__nor2_2 _13437_ (.A(_04320_),
    .B(_04321_),
    .Y(_04322_));
 sky130_fd_sc_hd__and2_1 _13438_ (.A(_04320_),
    .B(_04321_),
    .X(_04323_));
 sky130_fd_sc_hd__nor2_2 _13439_ (.A(_04322_),
    .B(_04323_),
    .Y(_04324_));
 sky130_fd_sc_hd__and2b_1 _13440_ (.A_N(_04187_),
    .B(_04324_),
    .X(_04326_));
 sky130_fd_sc_hd__inv_2 _13441_ (.A(_04326_),
    .Y(_04327_));
 sky130_fd_sc_hd__xnor2_2 _13442_ (.A(_04187_),
    .B(_04324_),
    .Y(_04328_));
 sky130_fd_sc_hd__and3_2 _13443_ (.A(_04316_),
    .B(_04317_),
    .C(_04328_),
    .X(_04329_));
 sky130_fd_sc_hd__inv_2 _13444_ (.A(_04329_),
    .Y(_04330_));
 sky130_fd_sc_hd__a21oi_4 _13445_ (.A1(_04316_),
    .A2(_04317_),
    .B1(_04328_),
    .Y(_04331_));
 sky130_fd_sc_hd__a211oi_4 _13446_ (.A1(_04192_),
    .A2(_04204_),
    .B1(_04329_),
    .C1(_04331_),
    .Y(_04332_));
 sky130_fd_sc_hd__o211a_2 _13447_ (.A1(_04329_),
    .A2(_04331_),
    .B1(_04192_),
    .C1(_04204_),
    .X(_04333_));
 sky130_fd_sc_hd__and2_4 _13448_ (.A(net392),
    .B(net699),
    .X(_04334_));
 sky130_fd_sc_hd__a22oi_1 _13449_ (.A1(net375),
    .A2(net715),
    .B1(net726),
    .B2(net366),
    .Y(_04335_));
 sky130_fd_sc_hd__and4_1 _13450_ (.A(net366),
    .B(net375),
    .C(net716),
    .D(net726),
    .X(_04337_));
 sky130_fd_sc_hd__nor2_1 _13451_ (.A(_04335_),
    .B(_04337_),
    .Y(_04338_));
 sky130_fd_sc_hd__a21oi_1 _13452_ (.A1(net384),
    .A2(net707),
    .B1(_04338_),
    .Y(_04339_));
 sky130_fd_sc_hd__and3_1 _13453_ (.A(net387),
    .B(net707),
    .C(_04338_),
    .X(_04340_));
 sky130_fd_sc_hd__nor2_1 _13454_ (.A(_04339_),
    .B(_04340_),
    .Y(_04341_));
 sky130_fd_sc_hd__or3_1 _13455_ (.A(_04210_),
    .B(_04213_),
    .C(_04341_),
    .X(_04342_));
 sky130_fd_sc_hd__o21ai_1 _13456_ (.A1(_04210_),
    .A2(_04213_),
    .B1(_04341_),
    .Y(_04343_));
 sky130_fd_sc_hd__and2_1 _13457_ (.A(_04342_),
    .B(_04343_),
    .X(_04344_));
 sky130_fd_sc_hd__nand2_1 _13458_ (.A(_04334_),
    .B(_04344_),
    .Y(_04345_));
 sky130_fd_sc_hd__or2_1 _13459_ (.A(_04334_),
    .B(_04344_),
    .X(_04346_));
 sky130_fd_sc_hd__nand2_1 _13460_ (.A(_04345_),
    .B(_04346_),
    .Y(_04348_));
 sky130_fd_sc_hd__a21oi_2 _13461_ (.A1(_04217_),
    .A2(_04219_),
    .B1(_04348_),
    .Y(_04349_));
 sky130_fd_sc_hd__and3_1 _13462_ (.A(_04217_),
    .B(_04219_),
    .C(_04348_),
    .X(_04350_));
 sky130_fd_sc_hd__nor2_2 _13463_ (.A(_04349_),
    .B(_04350_),
    .Y(_04351_));
 sky130_fd_sc_hd__nand2_1 _13464_ (.A(net400),
    .B(net689),
    .Y(_04352_));
 sky130_fd_sc_hd__xor2_2 _13465_ (.A(_04351_),
    .B(_04352_),
    .X(_04353_));
 sky130_fd_sc_hd__o21ba_1 _13466_ (.A1(_04195_),
    .A2(_04198_),
    .B1_N(_04196_),
    .X(_04354_));
 sky130_fd_sc_hd__a22oi_4 _13467_ (.A1(net351),
    .A2(net743),
    .B1(net752),
    .B2(net345),
    .Y(_04355_));
 sky130_fd_sc_hd__and4_1 _13468_ (.A(net345),
    .B(net351),
    .C(net743),
    .D(net752),
    .X(_04356_));
 sky130_fd_sc_hd__nor2_2 _13469_ (.A(_04355_),
    .B(_04356_),
    .Y(_04357_));
 sky130_fd_sc_hd__nand2_4 _13470_ (.A(net359),
    .B(net734),
    .Y(_04359_));
 sky130_fd_sc_hd__xnor2_4 _13471_ (.A(_04357_),
    .B(_04359_),
    .Y(_04360_));
 sky130_fd_sc_hd__and2b_1 _13472_ (.A_N(_04354_),
    .B(_04360_),
    .X(_04361_));
 sky130_fd_sc_hd__xnor2_2 _13473_ (.A(_04354_),
    .B(_04360_),
    .Y(_04362_));
 sky130_fd_sc_hd__o21ba_1 _13474_ (.A1(_04229_),
    .A2(_04232_),
    .B1_N(_04230_),
    .X(_04363_));
 sky130_fd_sc_hd__and2b_1 _13475_ (.A_N(_04363_),
    .B(_04362_),
    .X(_04364_));
 sky130_fd_sc_hd__xor2_1 _13476_ (.A(_04362_),
    .B(_04363_),
    .X(_04365_));
 sky130_fd_sc_hd__nor2_1 _13477_ (.A(_04234_),
    .B(_04237_),
    .Y(_04366_));
 sky130_fd_sc_hd__or2_2 _13478_ (.A(_04365_),
    .B(_04366_),
    .X(_04367_));
 sky130_fd_sc_hd__nand2_1 _13479_ (.A(_04365_),
    .B(_04366_),
    .Y(_04368_));
 sky130_fd_sc_hd__and2_1 _13480_ (.A(_04367_),
    .B(_04368_),
    .X(_04370_));
 sky130_fd_sc_hd__nand2_2 _13481_ (.A(_04241_),
    .B(_04370_),
    .Y(_04371_));
 sky130_fd_sc_hd__or2_1 _13482_ (.A(_04241_),
    .B(_04370_),
    .X(_04372_));
 sky130_fd_sc_hd__nand2_1 _13483_ (.A(_04371_),
    .B(_04372_),
    .Y(_04373_));
 sky130_fd_sc_hd__or2_4 _13484_ (.A(_04353_),
    .B(_04373_),
    .X(_04374_));
 sky130_fd_sc_hd__nand2_2 _13485_ (.A(_04353_),
    .B(_04373_),
    .Y(_04375_));
 sky130_fd_sc_hd__and3_4 _13486_ (.A(_04200_),
    .B(_04374_),
    .C(_04375_),
    .X(_04376_));
 sky130_fd_sc_hd__a21oi_4 _13487_ (.A1(_04374_),
    .A2(_04375_),
    .B1(_04200_),
    .Y(_04377_));
 sky130_fd_sc_hd__a211oi_4 _13488_ (.A1(_04244_),
    .A2(_04246_),
    .B1(_04376_),
    .C1(_04377_),
    .Y(_04378_));
 sky130_fd_sc_hd__o211a_2 _13489_ (.A1(_04376_),
    .A2(_04377_),
    .B1(_04244_),
    .C1(_04246_),
    .X(_04379_));
 sky130_fd_sc_hd__nor4_4 _13490_ (.A(_04332_),
    .B(_04333_),
    .C(_04378_),
    .D(_04379_),
    .Y(_04381_));
 sky130_fd_sc_hd__o22a_1 _13491_ (.A1(_04332_),
    .A2(_04333_),
    .B1(_04378_),
    .B2(_04379_),
    .X(_04382_));
 sky130_fd_sc_hd__nor2_1 _13492_ (.A(_04381_),
    .B(_04382_),
    .Y(_04383_));
 sky130_fd_sc_hd__o21a_2 _13493_ (.A1(_04207_),
    .A2(_04253_),
    .B1(_04383_),
    .X(_04384_));
 sky130_fd_sc_hd__nor3_1 _13494_ (.A(_04207_),
    .B(_04253_),
    .C(_04383_),
    .Y(_04385_));
 sky130_fd_sc_hd__nor2_2 _13495_ (.A(_04384_),
    .B(_04385_),
    .Y(_04386_));
 sky130_fd_sc_hd__nor2_2 _13496_ (.A(_04248_),
    .B(_04251_),
    .Y(_04387_));
 sky130_fd_sc_hd__and2b_2 _13497_ (.A_N(_04387_),
    .B(_04386_),
    .X(_04388_));
 sky130_fd_sc_hd__xnor2_2 _13498_ (.A(_04386_),
    .B(_04387_),
    .Y(_04389_));
 sky130_fd_sc_hd__o21a_1 _13499_ (.A1(_04255_),
    .A2(_04257_),
    .B1(_04389_),
    .X(_04390_));
 sky130_fd_sc_hd__nor3_2 _13500_ (.A(_04255_),
    .B(_04257_),
    .C(_04389_),
    .Y(_04392_));
 sky130_fd_sc_hd__nor2_1 _13501_ (.A(_04390_),
    .B(_04392_),
    .Y(_04393_));
 sky130_fd_sc_hd__o21ba_2 _13502_ (.A1(_04223_),
    .A2(_04225_),
    .B1_N(_04222_),
    .X(_04394_));
 sky130_fd_sc_hd__xnor2_2 _13503_ (.A(_04393_),
    .B(_04394_),
    .Y(_04395_));
 sky130_fd_sc_hd__or2_2 _13504_ (.A(_04259_),
    .B(_04262_),
    .X(_04396_));
 sky130_fd_sc_hd__nand2_4 _13505_ (.A(_04395_),
    .B(_04396_),
    .Y(_04397_));
 sky130_fd_sc_hd__or2_1 _13506_ (.A(_04395_),
    .B(_04396_),
    .X(_04398_));
 sky130_fd_sc_hd__nand2_2 _13507_ (.A(_04397_),
    .B(_04398_),
    .Y(_04399_));
 sky130_fd_sc_hd__and2b_1 _13508_ (.A_N(_04136_),
    .B(_04266_),
    .X(_04400_));
 sky130_fd_sc_hd__nor2_1 _13509_ (.A(_04135_),
    .B(_04264_),
    .Y(_04401_));
 sky130_fd_sc_hd__a211o_1 _13510_ (.A1(_04137_),
    .A2(_04400_),
    .B1(_04401_),
    .C1(_04265_),
    .X(_04403_));
 sky130_fd_sc_hd__and2_2 _13511_ (.A(_04138_),
    .B(_04400_),
    .X(_04404_));
 sky130_fd_sc_hd__a21oi_2 _13512_ (.A1(_03854_),
    .A2(_04404_),
    .B1(_04403_),
    .Y(_04405_));
 sky130_fd_sc_hd__nand2_1 _13513_ (.A(_04399_),
    .B(_04405_),
    .Y(_04406_));
 sky130_fd_sc_hd__or2_1 _13514_ (.A(_04399_),
    .B(_04405_),
    .X(_04407_));
 sky130_fd_sc_hd__a32o_1 _13515_ (.A1(net259),
    .A2(_04406_),
    .A3(_04407_),
    .B1(_04272_),
    .B2(_04275_),
    .X(_08655_));
 sky130_fd_sc_hd__mux2_8 _13516_ (.A0(_03350_),
    .A1(_03359_),
    .S(net567),
    .X(_04408_));
 sky130_fd_sc_hd__o21ai_1 _13517_ (.A1(net207),
    .A2(_04408_),
    .B1(net208),
    .Y(_04409_));
 sky130_fd_sc_hd__mux2_2 _13518_ (.A0(_03351_),
    .A1(_03354_),
    .S(net302),
    .X(_04410_));
 sky130_fd_sc_hd__nor2_1 _13519_ (.A(net306),
    .B(_04410_),
    .Y(_04411_));
 sky130_fd_sc_hd__a311o_1 _13520_ (.A1(net306),
    .A2(net570),
    .A3(_03353_),
    .B1(_04411_),
    .C1(net539),
    .X(_04413_));
 sky130_fd_sc_hd__a22o_1 _13521_ (.A1(net424),
    .A2(net656),
    .B1(net673),
    .B2(net408),
    .X(_04414_));
 sky130_fd_sc_hd__nand4_2 _13522_ (.A(net408),
    .B(net424),
    .C(net656),
    .D(net673),
    .Y(_04415_));
 sky130_fd_sc_hd__nand2_1 _13523_ (.A(net415),
    .B(net664),
    .Y(_04416_));
 sky130_fd_sc_hd__nand3b_1 _13524_ (.A_N(_04416_),
    .B(_04415_),
    .C(_04414_),
    .Y(_04417_));
 sky130_fd_sc_hd__a21bo_1 _13525_ (.A1(_04414_),
    .A2(_04415_),
    .B1_N(_04416_),
    .X(_04418_));
 sky130_fd_sc_hd__nand2_2 _13526_ (.A(_04277_),
    .B(_04279_),
    .Y(_04419_));
 sky130_fd_sc_hd__and3_1 _13527_ (.A(_04417_),
    .B(_04418_),
    .C(_04419_),
    .X(_04420_));
 sky130_fd_sc_hd__a21o_1 _13528_ (.A1(_04417_),
    .A2(_04418_),
    .B1(_04419_),
    .X(_04421_));
 sky130_fd_sc_hd__and2b_2 _13529_ (.A_N(_04420_),
    .B(_04421_),
    .X(_04422_));
 sky130_fd_sc_hd__a22oi_4 _13530_ (.A1(net445),
    .A2(net639),
    .B1(net648),
    .B2(net434),
    .Y(_04424_));
 sky130_fd_sc_hd__and4_2 _13531_ (.A(net434),
    .B(net445),
    .C(net639),
    .D(net648),
    .X(_04425_));
 sky130_fd_sc_hd__nor2_4 _13532_ (.A(_04424_),
    .B(_04425_),
    .Y(_04426_));
 sky130_fd_sc_hd__nand2_2 _13533_ (.A(net452),
    .B(net630),
    .Y(_04427_));
 sky130_fd_sc_hd__xnor2_4 _13534_ (.A(_04426_),
    .B(_04427_),
    .Y(_04428_));
 sky130_fd_sc_hd__xnor2_4 _13535_ (.A(_04422_),
    .B(_04428_),
    .Y(_04429_));
 sky130_fd_sc_hd__a21boi_4 _13536_ (.A1(_04284_),
    .A2(_04290_),
    .B1_N(_04283_),
    .Y(_04430_));
 sky130_fd_sc_hd__nor2_1 _13537_ (.A(_04429_),
    .B(_04430_),
    .Y(_04431_));
 sky130_fd_sc_hd__xnor2_4 _13538_ (.A(_04429_),
    .B(_04430_),
    .Y(_04432_));
 sky130_fd_sc_hd__a31o_1 _13539_ (.A1(net450),
    .A2(net636),
    .A3(_04288_),
    .B1(_04287_),
    .X(_04433_));
 sky130_fd_sc_hd__and3_1 _13540_ (.A(net459),
    .B(net619),
    .C(_04170_),
    .X(_04435_));
 sky130_fd_sc_hd__xor2_1 _13541_ (.A(_04433_),
    .B(_04435_),
    .X(_04436_));
 sky130_fd_sc_hd__clkinv_2 _13542_ (.A(_04436_),
    .Y(_04437_));
 sky130_fd_sc_hd__xnor2_4 _13543_ (.A(_04432_),
    .B(_04437_),
    .Y(_04438_));
 sky130_fd_sc_hd__a21oi_4 _13544_ (.A1(_04293_),
    .A2(_04307_),
    .B1(_04438_),
    .Y(_04439_));
 sky130_fd_sc_hd__and3_2 _13545_ (.A(_04293_),
    .B(_04307_),
    .C(_04438_),
    .X(_04440_));
 sky130_fd_sc_hd__a211oi_4 _13546_ (.A1(_04299_),
    .A2(_04302_),
    .B1(_04439_),
    .C1(_04440_),
    .Y(_04441_));
 sky130_fd_sc_hd__o211a_2 _13547_ (.A1(_04439_),
    .A2(_04440_),
    .B1(_04299_),
    .C1(_04302_),
    .X(_04442_));
 sky130_fd_sc_hd__a211o_4 _13548_ (.A1(_04309_),
    .A2(_04312_),
    .B1(_04441_),
    .C1(_04442_),
    .X(_04443_));
 sky130_fd_sc_hd__o211ai_4 _13549_ (.A1(_04441_),
    .A2(_04442_),
    .B1(_04309_),
    .C1(_04312_),
    .Y(_04444_));
 sky130_fd_sc_hd__a22oi_1 _13550_ (.A1(net333),
    .A2(net761),
    .B1(net773),
    .B2(net323),
    .Y(_04446_));
 sky130_fd_sc_hd__and4_1 _13551_ (.A(net323),
    .B(net333),
    .C(net765),
    .D(net776),
    .X(_04447_));
 sky130_fd_sc_hd__or2_1 _13552_ (.A(_04446_),
    .B(_04447_),
    .X(_04448_));
 sky130_fd_sc_hd__nand2_1 _13553_ (.A(net338),
    .B(net752),
    .Y(_04449_));
 sky130_fd_sc_hd__nor2_2 _13554_ (.A(_04448_),
    .B(_04449_),
    .Y(_04450_));
 sky130_fd_sc_hd__and2_1 _13555_ (.A(_04448_),
    .B(_04449_),
    .X(_04451_));
 sky130_fd_sc_hd__nor2_2 _13556_ (.A(_04450_),
    .B(_04451_),
    .Y(_04452_));
 sky130_fd_sc_hd__a21oi_4 _13557_ (.A1(_04443_),
    .A2(_04444_),
    .B1(_04452_),
    .Y(_04453_));
 sky130_fd_sc_hd__and3_2 _13558_ (.A(_04443_),
    .B(_04444_),
    .C(_04452_),
    .X(_04454_));
 sky130_fd_sc_hd__inv_2 _13559_ (.A(_04454_),
    .Y(_04455_));
 sky130_fd_sc_hd__a211oi_4 _13560_ (.A1(_04317_),
    .A2(_04330_),
    .B1(_04453_),
    .C1(_04454_),
    .Y(_04457_));
 sky130_fd_sc_hd__o211a_1 _13561_ (.A1(_04453_),
    .A2(_04454_),
    .B1(_04317_),
    .C1(_04330_),
    .X(_04458_));
 sky130_fd_sc_hd__nor2_4 _13562_ (.A(_04457_),
    .B(_04458_),
    .Y(_04459_));
 sky130_fd_sc_hd__a22oi_2 _13563_ (.A1(net375),
    .A2(net707),
    .B1(net716),
    .B2(net366),
    .Y(_04460_));
 sky130_fd_sc_hd__and4_2 _13564_ (.A(net366),
    .B(net375),
    .C(net707),
    .D(net716),
    .X(_04461_));
 sky130_fd_sc_hd__nor2_2 _13565_ (.A(_04460_),
    .B(_04461_),
    .Y(_04462_));
 sky130_fd_sc_hd__nand2_1 _13566_ (.A(net387),
    .B(net698),
    .Y(_04463_));
 sky130_fd_sc_hd__and3_1 _13567_ (.A(net387),
    .B(net698),
    .C(_04462_),
    .X(_04464_));
 sky130_fd_sc_hd__xnor2_2 _13568_ (.A(_04462_),
    .B(_04463_),
    .Y(_04465_));
 sky130_fd_sc_hd__or3_1 _13569_ (.A(_04337_),
    .B(_04340_),
    .C(_04465_),
    .X(_04466_));
 sky130_fd_sc_hd__o21ai_2 _13570_ (.A1(_04337_),
    .A2(_04340_),
    .B1(_04465_),
    .Y(_04468_));
 sky130_fd_sc_hd__and2_1 _13571_ (.A(_04466_),
    .B(_04468_),
    .X(_04469_));
 sky130_fd_sc_hd__nand3_2 _13572_ (.A(net392),
    .B(net690),
    .C(_04469_),
    .Y(_04470_));
 sky130_fd_sc_hd__a21o_1 _13573_ (.A1(net392),
    .A2(net690),
    .B1(_04469_),
    .X(_04471_));
 sky130_fd_sc_hd__nand2_1 _13574_ (.A(_04470_),
    .B(_04471_),
    .Y(_04472_));
 sky130_fd_sc_hd__a21oi_1 _13575_ (.A1(_04343_),
    .A2(_04345_),
    .B1(_04472_),
    .Y(_04473_));
 sky130_fd_sc_hd__and3_1 _13576_ (.A(_04343_),
    .B(_04345_),
    .C(_04472_),
    .X(_04474_));
 sky130_fd_sc_hd__nor2_1 _13577_ (.A(_04473_),
    .B(_04474_),
    .Y(_04475_));
 sky130_fd_sc_hd__nand2_1 _13578_ (.A(net400),
    .B(net680),
    .Y(_04476_));
 sky130_fd_sc_hd__xnor2_1 _13579_ (.A(_04475_),
    .B(_04476_),
    .Y(_04477_));
 sky130_fd_sc_hd__a22oi_2 _13580_ (.A1(net351),
    .A2(net734),
    .B1(net743),
    .B2(net345),
    .Y(_04479_));
 sky130_fd_sc_hd__and4_1 _13581_ (.A(net345),
    .B(net351),
    .C(net734),
    .D(net743),
    .X(_04480_));
 sky130_fd_sc_hd__nor2_1 _13582_ (.A(_04479_),
    .B(_04480_),
    .Y(_04481_));
 sky130_fd_sc_hd__nand2_2 _13583_ (.A(net362),
    .B(net726),
    .Y(_04482_));
 sky130_fd_sc_hd__xnor2_2 _13584_ (.A(_04481_),
    .B(_04482_),
    .Y(_04483_));
 sky130_fd_sc_hd__o21a_1 _13585_ (.A1(_04319_),
    .A2(_04322_),
    .B1(_04483_),
    .X(_04484_));
 sky130_fd_sc_hd__nor3_2 _13586_ (.A(_04319_),
    .B(_04322_),
    .C(_04483_),
    .Y(_04485_));
 sky130_fd_sc_hd__nor2_2 _13587_ (.A(_04484_),
    .B(_04485_),
    .Y(_04486_));
 sky130_fd_sc_hd__o21ba_2 _13588_ (.A1(_04355_),
    .A2(_04359_),
    .B1_N(_04356_),
    .X(_04487_));
 sky130_fd_sc_hd__xor2_4 _13589_ (.A(_04486_),
    .B(_04487_),
    .X(_04488_));
 sky130_fd_sc_hd__nor2_2 _13590_ (.A(_04361_),
    .B(_04364_),
    .Y(_04490_));
 sky130_fd_sc_hd__nor2_4 _13591_ (.A(_04488_),
    .B(_04490_),
    .Y(_04491_));
 sky130_fd_sc_hd__and2_1 _13592_ (.A(_04488_),
    .B(_04490_),
    .X(_04492_));
 sky130_fd_sc_hd__nor2_1 _13593_ (.A(_04491_),
    .B(_04492_),
    .Y(_04493_));
 sky130_fd_sc_hd__and2b_2 _13594_ (.A_N(_04367_),
    .B(_04493_),
    .X(_04494_));
 sky130_fd_sc_hd__xnor2_1 _13595_ (.A(_04367_),
    .B(_04493_),
    .Y(_04495_));
 sky130_fd_sc_hd__and2_2 _13596_ (.A(_04477_),
    .B(_04495_),
    .X(_04496_));
 sky130_fd_sc_hd__nor2_1 _13597_ (.A(_04477_),
    .B(_04495_),
    .Y(_04497_));
 sky130_fd_sc_hd__or2_1 _13598_ (.A(_04496_),
    .B(_04497_),
    .X(_04498_));
 sky130_fd_sc_hd__nor2_2 _13599_ (.A(_04327_),
    .B(_04498_),
    .Y(_04499_));
 sky130_fd_sc_hd__and2_1 _13600_ (.A(_04327_),
    .B(_04498_),
    .X(_04501_));
 sky130_fd_sc_hd__or2_2 _13601_ (.A(_04499_),
    .B(_04501_),
    .X(_04502_));
 sky130_fd_sc_hd__a21oi_4 _13602_ (.A1(_04371_),
    .A2(_04374_),
    .B1(_04502_),
    .Y(_04503_));
 sky130_fd_sc_hd__and3_1 _13603_ (.A(_04371_),
    .B(_04374_),
    .C(_04502_),
    .X(_04504_));
 sky130_fd_sc_hd__nor2_4 _13604_ (.A(_04503_),
    .B(_04504_),
    .Y(_04505_));
 sky130_fd_sc_hd__xor2_4 _13605_ (.A(_04459_),
    .B(_04505_),
    .X(_04506_));
 sky130_fd_sc_hd__o21ai_4 _13606_ (.A1(_04332_),
    .A2(_04381_),
    .B1(_04506_),
    .Y(_04507_));
 sky130_fd_sc_hd__or3_2 _13607_ (.A(_04332_),
    .B(_04381_),
    .C(_04506_),
    .X(_04508_));
 sky130_fd_sc_hd__o211ai_4 _13608_ (.A1(_04376_),
    .A2(_04378_),
    .B1(_04507_),
    .C1(_04508_),
    .Y(_04509_));
 sky130_fd_sc_hd__a211o_2 _13609_ (.A1(_04507_),
    .A2(_04508_),
    .B1(_04376_),
    .C1(_04378_),
    .X(_04510_));
 sky130_fd_sc_hd__o211a_2 _13610_ (.A1(_04384_),
    .A2(_04388_),
    .B1(_04509_),
    .C1(_04510_),
    .X(_04512_));
 sky130_fd_sc_hd__a211oi_4 _13611_ (.A1(_04509_),
    .A2(_04510_),
    .B1(_04384_),
    .C1(_04388_),
    .Y(_04513_));
 sky130_fd_sc_hd__nor2_4 _13612_ (.A(_04512_),
    .B(_04513_),
    .Y(_04514_));
 sky130_fd_sc_hd__a31o_4 _13613_ (.A1(net400),
    .A2(net689),
    .A3(_04351_),
    .B1(_04349_),
    .X(_04515_));
 sky130_fd_sc_hd__xor2_4 _13614_ (.A(_04514_),
    .B(_04515_),
    .X(_04516_));
 sky130_fd_sc_hd__o21ba_4 _13615_ (.A1(_04392_),
    .A2(_04394_),
    .B1_N(_04390_),
    .X(_04517_));
 sky130_fd_sc_hd__nand2b_1 _13616_ (.A_N(_04517_),
    .B(_04516_),
    .Y(_04518_));
 sky130_fd_sc_hd__and2b_1 _13617_ (.A_N(_04516_),
    .B(_04517_),
    .X(_04519_));
 sky130_fd_sc_hd__xnor2_4 _13618_ (.A(_04516_),
    .B(_04517_),
    .Y(_04520_));
 sky130_fd_sc_hd__nand2_1 _13619_ (.A(_04397_),
    .B(_04407_),
    .Y(_04521_));
 sky130_fd_sc_hd__nand2_1 _13620_ (.A(_04520_),
    .B(_04521_),
    .Y(_04523_));
 sky130_fd_sc_hd__or2_1 _13621_ (.A(_04520_),
    .B(_04521_),
    .X(_04524_));
 sky130_fd_sc_hd__a32o_1 _13622_ (.A1(net259),
    .A2(_04523_),
    .A3(_04524_),
    .B1(_04409_),
    .B2(_04413_),
    .X(_08656_));
 sky130_fd_sc_hd__mux2_1 _13623_ (.A0(_03523_),
    .A1(_03526_),
    .S(net568),
    .X(_04525_));
 sky130_fd_sc_hd__or2_2 _13624_ (.A(net553),
    .B(_04525_),
    .X(_04526_));
 sky130_fd_sc_hd__nor2_2 _13625_ (.A(net305),
    .B(_02642_),
    .Y(_04527_));
 sky130_fd_sc_hd__nand2_1 _13626_ (.A(net553),
    .B(_02641_),
    .Y(_04528_));
 sky130_fd_sc_hd__mux2_2 _13627_ (.A0(_03520_),
    .A1(_03522_),
    .S(net566),
    .X(_04529_));
 sky130_fd_sc_hd__nand2_1 _13628_ (.A(net568),
    .B(_03518_),
    .Y(_04530_));
 sky130_fd_sc_hd__o221a_1 _13629_ (.A1(_04528_),
    .A2(_04529_),
    .B1(_04530_),
    .B2(net207),
    .C1(net205),
    .X(_04531_));
 sky130_fd_sc_hd__a21oi_2 _13630_ (.A1(net538),
    .A2(_04526_),
    .B1(_04531_),
    .Y(_04533_));
 sky130_fd_sc_hd__a22oi_4 _13631_ (.A1(net424),
    .A2(net648),
    .B1(net664),
    .B2(net408),
    .Y(_04534_));
 sky130_fd_sc_hd__and4_4 _13632_ (.A(net408),
    .B(net424),
    .C(net648),
    .D(net664),
    .X(_04535_));
 sky130_fd_sc_hd__nand2_2 _13633_ (.A(net415),
    .B(net656),
    .Y(_04536_));
 sky130_fd_sc_hd__nor3_2 _13634_ (.A(_04534_),
    .B(_04535_),
    .C(_04536_),
    .Y(_04537_));
 sky130_fd_sc_hd__or3_2 _13635_ (.A(_04534_),
    .B(_04535_),
    .C(_04536_),
    .X(_04538_));
 sky130_fd_sc_hd__o21ai_2 _13636_ (.A1(_04534_),
    .A2(_04535_),
    .B1(_04536_),
    .Y(_04539_));
 sky130_fd_sc_hd__nand2_1 _13637_ (.A(_04415_),
    .B(_04417_),
    .Y(_04540_));
 sky130_fd_sc_hd__nand3_2 _13638_ (.A(_04538_),
    .B(_04539_),
    .C(_04540_),
    .Y(_04541_));
 sky130_fd_sc_hd__a21o_1 _13639_ (.A1(_04538_),
    .A2(_04539_),
    .B1(_04540_),
    .X(_04542_));
 sky130_fd_sc_hd__a22oi_2 _13640_ (.A1(net444),
    .A2(net630),
    .B1(net639),
    .B2(net434),
    .Y(_04544_));
 sky130_fd_sc_hd__and4_1 _13641_ (.A(net434),
    .B(net445),
    .C(net630),
    .D(net639),
    .X(_04545_));
 sky130_fd_sc_hd__nor2_1 _13642_ (.A(_04544_),
    .B(_04545_),
    .Y(_04546_));
 sky130_fd_sc_hd__nand2_2 _13643_ (.A(net452),
    .B(net623),
    .Y(_04547_));
 sky130_fd_sc_hd__xnor2_2 _13644_ (.A(_04546_),
    .B(_04547_),
    .Y(_04548_));
 sky130_fd_sc_hd__nand3_2 _13645_ (.A(_04541_),
    .B(_04542_),
    .C(_04548_),
    .Y(_04549_));
 sky130_fd_sc_hd__a21o_1 _13646_ (.A1(_04541_),
    .A2(_04542_),
    .B1(_04548_),
    .X(_04550_));
 sky130_fd_sc_hd__a21o_1 _13647_ (.A1(_04421_),
    .A2(_04428_),
    .B1(_04420_),
    .X(_04551_));
 sky130_fd_sc_hd__and3_1 _13648_ (.A(_04549_),
    .B(_04550_),
    .C(_04551_),
    .X(_04552_));
 sky130_fd_sc_hd__a21o_1 _13649_ (.A1(_04549_),
    .A2(_04550_),
    .B1(_04551_),
    .X(_04553_));
 sky130_fd_sc_hd__and2b_2 _13650_ (.A_N(_04552_),
    .B(_04553_),
    .X(_04555_));
 sky130_fd_sc_hd__a31o_4 _13651_ (.A1(net452),
    .A2(net630),
    .A3(_04426_),
    .B1(_04425_),
    .X(_04556_));
 sky130_fd_sc_hd__xnor2_4 _13652_ (.A(_04555_),
    .B(_04556_),
    .Y(_04557_));
 sky130_fd_sc_hd__o21bai_1 _13653_ (.A1(_04432_),
    .A2(_04437_),
    .B1_N(_04431_),
    .Y(_04558_));
 sky130_fd_sc_hd__and2b_1 _13654_ (.A_N(_04557_),
    .B(_04558_),
    .X(_04559_));
 sky130_fd_sc_hd__nand2b_1 _13655_ (.A_N(_04558_),
    .B(_04557_),
    .Y(_04560_));
 sky130_fd_sc_hd__nand2b_1 _13656_ (.A_N(_04559_),
    .B(_04560_),
    .Y(_04561_));
 sky130_fd_sc_hd__nand2b_1 _13657_ (.A_N(_04433_),
    .B(_04170_),
    .Y(_04562_));
 sky130_fd_sc_hd__and3_2 _13658_ (.A(net460),
    .B(net619),
    .C(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__xnor2_2 _13659_ (.A(_04561_),
    .B(_04563_),
    .Y(_04564_));
 sky130_fd_sc_hd__o21a_2 _13660_ (.A1(_04439_),
    .A2(_04441_),
    .B1(_04564_),
    .X(_04566_));
 sky130_fd_sc_hd__inv_2 _13661_ (.A(_04566_),
    .Y(_04567_));
 sky130_fd_sc_hd__or3_4 _13662_ (.A(_04439_),
    .B(_04441_),
    .C(_04564_),
    .X(_04568_));
 sky130_fd_sc_hd__a22oi_1 _13663_ (.A1(net333),
    .A2(net752),
    .B1(net765),
    .B2(net323),
    .Y(_04569_));
 sky130_fd_sc_hd__and4_1 _13664_ (.A(net323),
    .B(net333),
    .C(net752),
    .D(net765),
    .X(_04570_));
 sky130_fd_sc_hd__or2_1 _13665_ (.A(_04569_),
    .B(_04570_),
    .X(_04571_));
 sky130_fd_sc_hd__nand2_1 _13666_ (.A(net338),
    .B(net743),
    .Y(_04572_));
 sky130_fd_sc_hd__nor2_2 _13667_ (.A(_04571_),
    .B(_04572_),
    .Y(_04573_));
 sky130_fd_sc_hd__and2_1 _13668_ (.A(_04571_),
    .B(_04572_),
    .X(_04574_));
 sky130_fd_sc_hd__nor2_2 _13669_ (.A(_04573_),
    .B(_04574_),
    .Y(_04575_));
 sky130_fd_sc_hd__a21oi_4 _13670_ (.A1(_04567_),
    .A2(_04568_),
    .B1(_04575_),
    .Y(_04577_));
 sky130_fd_sc_hd__and3_4 _13671_ (.A(_04567_),
    .B(_04568_),
    .C(_04575_),
    .X(_04578_));
 sky130_fd_sc_hd__a211oi_4 _13672_ (.A1(_04443_),
    .A2(_04455_),
    .B1(_04577_),
    .C1(_04578_),
    .Y(_04579_));
 sky130_fd_sc_hd__o211a_1 _13673_ (.A1(_04577_),
    .A2(_04578_),
    .B1(_04443_),
    .C1(_04455_),
    .X(_04580_));
 sky130_fd_sc_hd__a22oi_2 _13674_ (.A1(net351),
    .A2(net726),
    .B1(net734),
    .B2(net346),
    .Y(_04581_));
 sky130_fd_sc_hd__and4_1 _13675_ (.A(net346),
    .B(net351),
    .C(net726),
    .D(net734),
    .X(_04582_));
 sky130_fd_sc_hd__nor2_1 _13676_ (.A(_04581_),
    .B(_04582_),
    .Y(_04583_));
 sky130_fd_sc_hd__nand2_1 _13677_ (.A(net362),
    .B(net716),
    .Y(_04584_));
 sky130_fd_sc_hd__xnor2_1 _13678_ (.A(_04583_),
    .B(_04584_),
    .Y(_04585_));
 sky130_fd_sc_hd__o21a_1 _13679_ (.A1(_04447_),
    .A2(_04450_),
    .B1(_04585_),
    .X(_04586_));
 sky130_fd_sc_hd__nor3_1 _13680_ (.A(_04447_),
    .B(_04450_),
    .C(_04585_),
    .Y(_04588_));
 sky130_fd_sc_hd__nor2_1 _13681_ (.A(_04586_),
    .B(_04588_),
    .Y(_04589_));
 sky130_fd_sc_hd__o21ba_1 _13682_ (.A1(_04479_),
    .A2(_04482_),
    .B1_N(_04480_),
    .X(_04590_));
 sky130_fd_sc_hd__xor2_1 _13683_ (.A(_04589_),
    .B(_04590_),
    .X(_04591_));
 sky130_fd_sc_hd__o21ba_1 _13684_ (.A1(_04485_),
    .A2(_04487_),
    .B1_N(_04484_),
    .X(_04592_));
 sky130_fd_sc_hd__or2_2 _13685_ (.A(_04591_),
    .B(_04592_),
    .X(_04593_));
 sky130_fd_sc_hd__nand2_1 _13686_ (.A(_04591_),
    .B(_04592_),
    .Y(_04594_));
 sky130_fd_sc_hd__and2_2 _13687_ (.A(_04593_),
    .B(_04594_),
    .X(_04595_));
 sky130_fd_sc_hd__xor2_2 _13688_ (.A(_04491_),
    .B(_04595_),
    .X(_04596_));
 sky130_fd_sc_hd__nand2_8 _13689_ (.A(net384),
    .B(net686),
    .Y(_04597_));
 sky130_fd_sc_hd__a22oi_4 _13690_ (.A1(net376),
    .A2(net698),
    .B1(net708),
    .B2(net367),
    .Y(_04599_));
 sky130_fd_sc_hd__and4_2 _13691_ (.A(net367),
    .B(net376),
    .C(net698),
    .D(net708),
    .X(_04600_));
 sky130_fd_sc_hd__o21a_1 _13692_ (.A1(_04599_),
    .A2(_04600_),
    .B1(_04597_),
    .X(_04601_));
 sky130_fd_sc_hd__nor3_2 _13693_ (.A(_04597_),
    .B(_04599_),
    .C(_04600_),
    .Y(_04602_));
 sky130_fd_sc_hd__nor2_1 _13694_ (.A(_04601_),
    .B(_04602_),
    .Y(_04603_));
 sky130_fd_sc_hd__or3_1 _13695_ (.A(_04461_),
    .B(_04464_),
    .C(_04603_),
    .X(_04604_));
 sky130_fd_sc_hd__o21ai_2 _13696_ (.A1(_04461_),
    .A2(_04464_),
    .B1(_04603_),
    .Y(_04605_));
 sky130_fd_sc_hd__and2_1 _13697_ (.A(_04604_),
    .B(_04605_),
    .X(_04606_));
 sky130_fd_sc_hd__nand3_2 _13698_ (.A(net392),
    .B(net683),
    .C(_04606_),
    .Y(_04607_));
 sky130_fd_sc_hd__a21o_1 _13699_ (.A1(net392),
    .A2(net683),
    .B1(_04606_),
    .X(_04608_));
 sky130_fd_sc_hd__nand2_1 _13700_ (.A(_04607_),
    .B(_04608_),
    .Y(_04610_));
 sky130_fd_sc_hd__a21oi_2 _13701_ (.A1(_04468_),
    .A2(_04470_),
    .B1(_04610_),
    .Y(_04611_));
 sky130_fd_sc_hd__and3_1 _13702_ (.A(_04468_),
    .B(_04470_),
    .C(_04610_),
    .X(_04612_));
 sky130_fd_sc_hd__nor2_2 _13703_ (.A(_04611_),
    .B(_04612_),
    .Y(_04613_));
 sky130_fd_sc_hd__nand2_1 _13704_ (.A(net400),
    .B(net670),
    .Y(_04614_));
 sky130_fd_sc_hd__xnor2_1 _13705_ (.A(_04613_),
    .B(_04614_),
    .Y(_04615_));
 sky130_fd_sc_hd__nand2_2 _13706_ (.A(_04596_),
    .B(_04615_),
    .Y(_04616_));
 sky130_fd_sc_hd__or2_2 _13707_ (.A(_04596_),
    .B(_04615_),
    .X(_04617_));
 sky130_fd_sc_hd__o211a_4 _13708_ (.A1(_04494_),
    .A2(_04496_),
    .B1(_04616_),
    .C1(_04617_),
    .X(_04618_));
 sky130_fd_sc_hd__a211oi_4 _13709_ (.A1(_04616_),
    .A2(_04617_),
    .B1(_04494_),
    .C1(_04496_),
    .Y(_04619_));
 sky130_fd_sc_hd__nor4_2 _13710_ (.A(_04579_),
    .B(_04580_),
    .C(_04618_),
    .D(_04619_),
    .Y(_04621_));
 sky130_fd_sc_hd__o22a_2 _13711_ (.A1(_04579_),
    .A2(_04580_),
    .B1(_04618_),
    .B2(_04619_),
    .X(_04622_));
 sky130_fd_sc_hd__a21oi_4 _13712_ (.A1(_04459_),
    .A2(_04505_),
    .B1(_04457_),
    .Y(_04623_));
 sky130_fd_sc_hd__or3_4 _13713_ (.A(net117),
    .B(_04622_),
    .C(_04623_),
    .X(_04624_));
 sky130_fd_sc_hd__o21ai_4 _13714_ (.A1(net117),
    .A2(_04622_),
    .B1(_04623_),
    .Y(_04625_));
 sky130_fd_sc_hd__o211ai_4 _13715_ (.A1(_04499_),
    .A2(_04503_),
    .B1(_04624_),
    .C1(_04625_),
    .Y(_04626_));
 sky130_fd_sc_hd__a211o_1 _13716_ (.A1(_04624_),
    .A2(_04625_),
    .B1(_04499_),
    .C1(_04503_),
    .X(_04627_));
 sky130_fd_sc_hd__and2_2 _13717_ (.A(_04626_),
    .B(_04627_),
    .X(_04628_));
 sky130_fd_sc_hd__nand2_2 _13718_ (.A(_04507_),
    .B(_04509_),
    .Y(_04629_));
 sky130_fd_sc_hd__nand2_1 _13719_ (.A(_04628_),
    .B(_04629_),
    .Y(_04630_));
 sky130_fd_sc_hd__xnor2_2 _13720_ (.A(_04628_),
    .B(_04629_),
    .Y(_04632_));
 sky130_fd_sc_hd__o21ba_2 _13721_ (.A1(_04474_),
    .A2(_04476_),
    .B1_N(_04473_),
    .X(_04633_));
 sky130_fd_sc_hd__or2_1 _13722_ (.A(_04632_),
    .B(_04633_),
    .X(_04634_));
 sky130_fd_sc_hd__xnor2_2 _13723_ (.A(_04632_),
    .B(_04633_),
    .Y(_04635_));
 sky130_fd_sc_hd__a21oi_2 _13724_ (.A1(_04514_),
    .A2(_04515_),
    .B1(_04512_),
    .Y(_04636_));
 sky130_fd_sc_hd__nor2_2 _13725_ (.A(_04635_),
    .B(_04636_),
    .Y(_04637_));
 sky130_fd_sc_hd__and2_1 _13726_ (.A(_04635_),
    .B(_04636_),
    .X(_04638_));
 sky130_fd_sc_hd__or2_2 _13727_ (.A(_04637_),
    .B(_04638_),
    .X(_04639_));
 sky130_fd_sc_hd__a21oi_2 _13728_ (.A1(_04397_),
    .A2(_04518_),
    .B1(_04519_),
    .Y(_04640_));
 sky130_fd_sc_hd__nand2b_2 _13729_ (.A_N(_04399_),
    .B(_04520_),
    .Y(_04641_));
 sky130_fd_sc_hd__o21ba_1 _13730_ (.A1(_04405_),
    .A2(_04641_),
    .B1_N(_04640_),
    .X(_04643_));
 sky130_fd_sc_hd__nand2_1 _13731_ (.A(_04639_),
    .B(_04643_),
    .Y(_04644_));
 sky130_fd_sc_hd__or2_1 _13732_ (.A(_04639_),
    .B(_04643_),
    .X(_04645_));
 sky130_fd_sc_hd__a31o_1 _13733_ (.A1(net259),
    .A2(_04644_),
    .A3(_04645_),
    .B1(_04533_),
    .X(_08657_));
 sky130_fd_sc_hd__a22oi_2 _13734_ (.A1(net424),
    .A2(net640),
    .B1(net656),
    .B2(net408),
    .Y(_04646_));
 sky130_fd_sc_hd__and4_2 _13735_ (.A(net408),
    .B(net424),
    .C(net640),
    .D(net656),
    .X(_04647_));
 sky130_fd_sc_hd__nor2_2 _13736_ (.A(_04646_),
    .B(_04647_),
    .Y(_04648_));
 sky130_fd_sc_hd__nand2_1 _13737_ (.A(net415),
    .B(net648),
    .Y(_04649_));
 sky130_fd_sc_hd__and3_1 _13738_ (.A(net415),
    .B(net648),
    .C(_04648_),
    .X(_04650_));
 sky130_fd_sc_hd__xnor2_2 _13739_ (.A(_04648_),
    .B(_04649_),
    .Y(_04651_));
 sky130_fd_sc_hd__o21a_2 _13740_ (.A1(_04535_),
    .A2(_04537_),
    .B1(_04651_),
    .X(_04653_));
 sky130_fd_sc_hd__nor3_2 _13741_ (.A(_04535_),
    .B(_04537_),
    .C(_04651_),
    .Y(_04654_));
 sky130_fd_sc_hd__nor2_4 _13742_ (.A(_04653_),
    .B(_04654_),
    .Y(_04655_));
 sky130_fd_sc_hd__a22oi_1 _13743_ (.A1(net444),
    .A2(net623),
    .B1(net630),
    .B2(net434),
    .Y(_04656_));
 sky130_fd_sc_hd__nand2_1 _13744_ (.A(net434),
    .B(net622),
    .Y(_04657_));
 sky130_fd_sc_hd__and4_1 _13745_ (.A(net435),
    .B(net445),
    .C(net623),
    .D(net630),
    .X(_04658_));
 sky130_fd_sc_hd__or2_1 _13746_ (.A(_04656_),
    .B(_04658_),
    .X(_04659_));
 sky130_fd_sc_hd__clkinv_2 _13747_ (.A(_04659_),
    .Y(_04660_));
 sky130_fd_sc_hd__xnor2_4 _13748_ (.A(_04655_),
    .B(_04660_),
    .Y(_04661_));
 sky130_fd_sc_hd__nand2_1 _13749_ (.A(_04541_),
    .B(_04549_),
    .Y(_04662_));
 sky130_fd_sc_hd__a21o_1 _13750_ (.A1(_04541_),
    .A2(_04549_),
    .B1(_04661_),
    .X(_04664_));
 sky130_fd_sc_hd__xnor2_2 _13751_ (.A(_04661_),
    .B(_04662_),
    .Y(_04665_));
 sky130_fd_sc_hd__o21ba_1 _13752_ (.A1(_04544_),
    .A2(_04547_),
    .B1_N(_04545_),
    .X(_04666_));
 sky130_fd_sc_hd__nand2b_1 _13753_ (.A_N(_04666_),
    .B(_04665_),
    .Y(_04667_));
 sky130_fd_sc_hd__xnor2_1 _13754_ (.A(_04665_),
    .B(_04666_),
    .Y(_04668_));
 sky130_fd_sc_hd__a21oi_1 _13755_ (.A1(_04553_),
    .A2(_04556_),
    .B1(_04552_),
    .Y(_04669_));
 sky130_fd_sc_hd__and2b_1 _13756_ (.A_N(_04669_),
    .B(_04668_),
    .X(_04670_));
 sky130_fd_sc_hd__and2b_1 _13757_ (.A_N(_04668_),
    .B(_04669_),
    .X(_04671_));
 sky130_fd_sc_hd__or2_4 _13758_ (.A(_04670_),
    .B(_04671_),
    .X(_04672_));
 sky130_fd_sc_hd__a21oi_2 _13759_ (.A1(_04560_),
    .A2(_04563_),
    .B1(_04559_),
    .Y(_04673_));
 sky130_fd_sc_hd__nor2_2 _13760_ (.A(_04672_),
    .B(_04673_),
    .Y(_04675_));
 sky130_fd_sc_hd__and2_1 _13761_ (.A(_04672_),
    .B(_04673_),
    .X(_04676_));
 sky130_fd_sc_hd__nor2_4 _13762_ (.A(_04675_),
    .B(_04676_),
    .Y(_04677_));
 sky130_fd_sc_hd__a22oi_4 _13763_ (.A1(net333),
    .A2(net743),
    .B1(net751),
    .B2(net323),
    .Y(_04678_));
 sky130_fd_sc_hd__and4_1 _13764_ (.A(net323),
    .B(net333),
    .C(net742),
    .D(net751),
    .X(_04679_));
 sky130_fd_sc_hd__nor2_2 _13765_ (.A(_04678_),
    .B(_04679_),
    .Y(_04680_));
 sky130_fd_sc_hd__nand2_4 _13766_ (.A(net338),
    .B(net734),
    .Y(_04681_));
 sky130_fd_sc_hd__xnor2_4 _13767_ (.A(_04680_),
    .B(_04681_),
    .Y(_04682_));
 sky130_fd_sc_hd__xor2_4 _13768_ (.A(_04677_),
    .B(_04682_),
    .X(_04683_));
 sky130_fd_sc_hd__o21ai_2 _13769_ (.A1(_04566_),
    .A2(_04578_),
    .B1(_04683_),
    .Y(_04684_));
 sky130_fd_sc_hd__or3_1 _13770_ (.A(_04566_),
    .B(_04578_),
    .C(_04683_),
    .X(_04686_));
 sky130_fd_sc_hd__nand2_2 _13771_ (.A(_04684_),
    .B(_04686_),
    .Y(_04687_));
 sky130_fd_sc_hd__a22oi_2 _13772_ (.A1(net351),
    .A2(net716),
    .B1(net726),
    .B2(net345),
    .Y(_04688_));
 sky130_fd_sc_hd__and4_1 _13773_ (.A(net345),
    .B(net351),
    .C(net716),
    .D(net726),
    .X(_04689_));
 sky130_fd_sc_hd__nor2_1 _13774_ (.A(_04688_),
    .B(_04689_),
    .Y(_04690_));
 sky130_fd_sc_hd__nand2_1 _13775_ (.A(net359),
    .B(net707),
    .Y(_04691_));
 sky130_fd_sc_hd__xnor2_1 _13776_ (.A(_04690_),
    .B(_04691_),
    .Y(_04692_));
 sky130_fd_sc_hd__o21a_1 _13777_ (.A1(_04570_),
    .A2(_04573_),
    .B1(_04692_),
    .X(_04693_));
 sky130_fd_sc_hd__nor3_1 _13778_ (.A(_04570_),
    .B(_04573_),
    .C(_04692_),
    .Y(_04694_));
 sky130_fd_sc_hd__nor2_1 _13779_ (.A(_04693_),
    .B(_04694_),
    .Y(_04695_));
 sky130_fd_sc_hd__o21ba_1 _13780_ (.A1(_04581_),
    .A2(_04584_),
    .B1_N(_04582_),
    .X(_04697_));
 sky130_fd_sc_hd__xor2_1 _13781_ (.A(_04695_),
    .B(_04697_),
    .X(_04698_));
 sky130_fd_sc_hd__o21ba_1 _13782_ (.A1(_04588_),
    .A2(_04590_),
    .B1_N(_04586_),
    .X(_04699_));
 sky130_fd_sc_hd__nor2_1 _13783_ (.A(_04698_),
    .B(_04699_),
    .Y(_04700_));
 sky130_fd_sc_hd__and2_1 _13784_ (.A(_04698_),
    .B(_04699_),
    .X(_04701_));
 sky130_fd_sc_hd__nor2_1 _13785_ (.A(_04700_),
    .B(_04701_),
    .Y(_04702_));
 sky130_fd_sc_hd__and2b_1 _13786_ (.A_N(_04593_),
    .B(_04702_),
    .X(_04703_));
 sky130_fd_sc_hd__xnor2_1 _13787_ (.A(_04593_),
    .B(_04702_),
    .Y(_04704_));
 sky130_fd_sc_hd__a22oi_2 _13788_ (.A1(net380),
    .A2(net690),
    .B1(net698),
    .B2(net371),
    .Y(_04705_));
 sky130_fd_sc_hd__and4_1 _13789_ (.A(net371),
    .B(net380),
    .C(net690),
    .D(net700),
    .X(_04706_));
 sky130_fd_sc_hd__nor2_1 _13790_ (.A(_04705_),
    .B(_04706_),
    .Y(_04708_));
 sky130_fd_sc_hd__nand2_1 _13791_ (.A(net387),
    .B(net680),
    .Y(_04709_));
 sky130_fd_sc_hd__xnor2_1 _13792_ (.A(_04708_),
    .B(_04709_),
    .Y(_04710_));
 sky130_fd_sc_hd__or3_1 _13793_ (.A(_04600_),
    .B(_04602_),
    .C(_04710_),
    .X(_04711_));
 sky130_fd_sc_hd__o21ai_2 _13794_ (.A1(_04600_),
    .A2(_04602_),
    .B1(_04710_),
    .Y(_04712_));
 sky130_fd_sc_hd__and2_1 _13795_ (.A(_04711_),
    .B(_04712_),
    .X(_04713_));
 sky130_fd_sc_hd__nand3_2 _13796_ (.A(net393),
    .B(net670),
    .C(_04713_),
    .Y(_04714_));
 sky130_fd_sc_hd__a21o_1 _13797_ (.A1(net393),
    .A2(net670),
    .B1(_04713_),
    .X(_04715_));
 sky130_fd_sc_hd__nand2_1 _13798_ (.A(_04714_),
    .B(_04715_),
    .Y(_04716_));
 sky130_fd_sc_hd__a21oi_2 _13799_ (.A1(_04605_),
    .A2(_04607_),
    .B1(_04716_),
    .Y(_04717_));
 sky130_fd_sc_hd__and3_1 _13800_ (.A(_04605_),
    .B(_04607_),
    .C(_04716_),
    .X(_04719_));
 sky130_fd_sc_hd__nor2_2 _13801_ (.A(_04717_),
    .B(_04719_),
    .Y(_04720_));
 sky130_fd_sc_hd__nand2_1 _13802_ (.A(net401),
    .B(net662),
    .Y(_04721_));
 sky130_fd_sc_hd__xnor2_1 _13803_ (.A(_04720_),
    .B(_04721_),
    .Y(_04722_));
 sky130_fd_sc_hd__and2_1 _13804_ (.A(_04704_),
    .B(_04722_),
    .X(_04723_));
 sky130_fd_sc_hd__nor2_1 _13805_ (.A(_04704_),
    .B(_04722_),
    .Y(_04724_));
 sky130_fd_sc_hd__or2_2 _13806_ (.A(_04723_),
    .B(_04724_),
    .X(_04725_));
 sky130_fd_sc_hd__a21boi_4 _13807_ (.A1(_04491_),
    .A2(_04595_),
    .B1_N(_04616_),
    .Y(_04726_));
 sky130_fd_sc_hd__nor2_2 _13808_ (.A(_04725_),
    .B(_04726_),
    .Y(_04727_));
 sky130_fd_sc_hd__and2_1 _13809_ (.A(_04725_),
    .B(_04726_),
    .X(_04728_));
 sky130_fd_sc_hd__or2_2 _13810_ (.A(_04727_),
    .B(_04728_),
    .X(_04730_));
 sky130_fd_sc_hd__or2_1 _13811_ (.A(_04687_),
    .B(_04730_),
    .X(_04731_));
 sky130_fd_sc_hd__xor2_2 _13812_ (.A(_04687_),
    .B(_04730_),
    .X(_04732_));
 sky130_fd_sc_hd__o21ai_2 _13813_ (.A1(_04579_),
    .A2(_04621_),
    .B1(_04732_),
    .Y(_04733_));
 sky130_fd_sc_hd__or3_1 _13814_ (.A(_04579_),
    .B(_04621_),
    .C(_04732_),
    .X(_04734_));
 sky130_fd_sc_hd__and2_2 _13815_ (.A(_04733_),
    .B(_04734_),
    .X(_04735_));
 sky130_fd_sc_hd__nand2_1 _13816_ (.A(_04618_),
    .B(_04735_),
    .Y(_04736_));
 sky130_fd_sc_hd__xnor2_4 _13817_ (.A(_04618_),
    .B(_04735_),
    .Y(_04737_));
 sky130_fd_sc_hd__nand2_4 _13818_ (.A(_04624_),
    .B(_04626_),
    .Y(_04738_));
 sky130_fd_sc_hd__and2b_1 _13819_ (.A_N(_04737_),
    .B(_04738_),
    .X(_04739_));
 sky130_fd_sc_hd__xor2_4 _13820_ (.A(_04737_),
    .B(_04738_),
    .X(_04741_));
 sky130_fd_sc_hd__a31o_4 _13821_ (.A1(net400),
    .A2(net670),
    .A3(_04613_),
    .B1(_04611_),
    .X(_04742_));
 sky130_fd_sc_hd__and2b_1 _13822_ (.A_N(_04741_),
    .B(_04742_),
    .X(_04743_));
 sky130_fd_sc_hd__xor2_4 _13823_ (.A(_04741_),
    .B(_04742_),
    .X(_04744_));
 sky130_fd_sc_hd__nand2_2 _13824_ (.A(_04630_),
    .B(_04634_),
    .Y(_04745_));
 sky130_fd_sc_hd__nand2b_1 _13825_ (.A_N(_04745_),
    .B(_04744_),
    .Y(_04746_));
 sky130_fd_sc_hd__a21oi_1 _13826_ (.A1(_04630_),
    .A2(_04634_),
    .B1(_04744_),
    .Y(_04747_));
 sky130_fd_sc_hd__xor2_4 _13827_ (.A(_04744_),
    .B(_04745_),
    .X(_04748_));
 sky130_fd_sc_hd__and2b_1 _13828_ (.A_N(_04637_),
    .B(_04645_),
    .X(_04749_));
 sky130_fd_sc_hd__nand2_1 _13829_ (.A(_04748_),
    .B(_04749_),
    .Y(_04750_));
 sky130_fd_sc_hd__or2_1 _13830_ (.A(_04748_),
    .B(_04749_),
    .X(_04752_));
 sky130_fd_sc_hd__mux2_1 _13831_ (.A0(_03675_),
    .A1(_03683_),
    .S(net570),
    .X(_04753_));
 sky130_fd_sc_hd__nor2_1 _13832_ (.A(net553),
    .B(_04753_),
    .Y(_04754_));
 sky130_fd_sc_hd__mux2_2 _13833_ (.A0(_03676_),
    .A1(_03679_),
    .S(net300),
    .X(_04755_));
 sky130_fd_sc_hd__inv_2 _13834_ (.A(_04755_),
    .Y(_04756_));
 sky130_fd_sc_hd__a32o_1 _13835_ (.A1(net553),
    .A2(_02643_),
    .A3(_04756_),
    .B1(_04754_),
    .B2(_03685_),
    .X(_04757_));
 sky130_fd_sc_hd__a31o_1 _13836_ (.A1(net259),
    .A2(_04750_),
    .A3(_04752_),
    .B1(_04757_),
    .X(_08658_));
 sky130_fd_sc_hd__or3_2 _13837_ (.A(net568),
    .B(net585),
    .C(_03190_),
    .X(_04758_));
 sky130_fd_sc_hd__mux2_1 _13838_ (.A0(_03688_),
    .A1(_03693_),
    .S(net301),
    .X(_04759_));
 sky130_fd_sc_hd__mux2_2 _13839_ (.A0(_04758_),
    .A1(_04759_),
    .S(net308),
    .X(_04760_));
 sky130_fd_sc_hd__mux2_1 _13840_ (.A0(_03694_),
    .A1(_03697_),
    .S(net300),
    .X(_04762_));
 sky130_fd_sc_hd__or2_1 _13841_ (.A(net204),
    .B(_04762_),
    .X(_04763_));
 sky130_fd_sc_hd__a22o_2 _13842_ (.A1(net537),
    .A2(_04760_),
    .B1(_04763_),
    .B2(net205),
    .X(_04764_));
 sky130_fd_sc_hd__a22oi_1 _13843_ (.A1(net424),
    .A2(net630),
    .B1(net649),
    .B2(net408),
    .Y(_04765_));
 sky130_fd_sc_hd__and4_1 _13844_ (.A(net408),
    .B(net424),
    .C(net630),
    .D(net649),
    .X(_04766_));
 sky130_fd_sc_hd__nor2_1 _13845_ (.A(_04765_),
    .B(_04766_),
    .Y(_04767_));
 sky130_fd_sc_hd__nand2_1 _13846_ (.A(net415),
    .B(net639),
    .Y(_04768_));
 sky130_fd_sc_hd__and3_1 _13847_ (.A(net415),
    .B(net639),
    .C(_04767_),
    .X(_04769_));
 sky130_fd_sc_hd__xnor2_1 _13848_ (.A(_04767_),
    .B(_04768_),
    .Y(_04770_));
 sky130_fd_sc_hd__nor3_1 _13849_ (.A(_04647_),
    .B(_04650_),
    .C(_04770_),
    .Y(_04771_));
 sky130_fd_sc_hd__o21a_2 _13850_ (.A1(_04647_),
    .A2(_04650_),
    .B1(_04770_),
    .X(_04773_));
 sky130_fd_sc_hd__nor2_2 _13851_ (.A(_04771_),
    .B(_04773_),
    .Y(_04774_));
 sky130_fd_sc_hd__and3_1 _13852_ (.A(net434),
    .B(net623),
    .C(_04774_),
    .X(_04775_));
 sky130_fd_sc_hd__xor2_2 _13853_ (.A(_04657_),
    .B(_04774_),
    .X(_04776_));
 sky130_fd_sc_hd__a21o_1 _13854_ (.A1(_04655_),
    .A2(_04660_),
    .B1(_04653_),
    .X(_04777_));
 sky130_fd_sc_hd__and2b_1 _13855_ (.A_N(_04776_),
    .B(_04777_),
    .X(_04778_));
 sky130_fd_sc_hd__xnor2_1 _13856_ (.A(_04776_),
    .B(_04777_),
    .Y(_04779_));
 sky130_fd_sc_hd__and2_1 _13857_ (.A(_04658_),
    .B(_04779_),
    .X(_04780_));
 sky130_fd_sc_hd__nor2_1 _13858_ (.A(_04658_),
    .B(_04779_),
    .Y(_04781_));
 sky130_fd_sc_hd__or2_1 _13859_ (.A(_04780_),
    .B(_04781_),
    .X(_04782_));
 sky130_fd_sc_hd__a21o_2 _13860_ (.A1(_04664_),
    .A2(_04667_),
    .B1(_04782_),
    .X(_04784_));
 sky130_fd_sc_hd__nand3_1 _13861_ (.A(_04664_),
    .B(_04667_),
    .C(_04782_),
    .Y(_04785_));
 sky130_fd_sc_hd__and3_4 _13862_ (.A(_04670_),
    .B(_04784_),
    .C(_04785_),
    .X(_04786_));
 sky130_fd_sc_hd__a21o_2 _13863_ (.A1(_04784_),
    .A2(_04785_),
    .B1(_04670_),
    .X(_04787_));
 sky130_fd_sc_hd__nand2b_1 _13864_ (.A_N(_04786_),
    .B(_04787_),
    .Y(_04788_));
 sky130_fd_sc_hd__a22oi_4 _13865_ (.A1(net331),
    .A2(net734),
    .B1(net743),
    .B2(net321),
    .Y(_04789_));
 sky130_fd_sc_hd__and4_1 _13866_ (.A(net321),
    .B(net331),
    .C(net734),
    .D(net743),
    .X(_04790_));
 sky130_fd_sc_hd__nor2_2 _13867_ (.A(_04789_),
    .B(_04790_),
    .Y(_04791_));
 sky130_fd_sc_hd__nand2_4 _13868_ (.A(net338),
    .B(net726),
    .Y(_04792_));
 sky130_fd_sc_hd__xnor2_4 _13869_ (.A(_04791_),
    .B(_04792_),
    .Y(_04793_));
 sky130_fd_sc_hd__xnor2_1 _13870_ (.A(_04788_),
    .B(_04793_),
    .Y(_04795_));
 sky130_fd_sc_hd__a21o_1 _13871_ (.A1(_04677_),
    .A2(_04682_),
    .B1(_04675_),
    .X(_04796_));
 sky130_fd_sc_hd__nand2_1 _13872_ (.A(_04795_),
    .B(_04796_),
    .Y(_04797_));
 sky130_fd_sc_hd__or2_1 _13873_ (.A(_04795_),
    .B(_04796_),
    .X(_04798_));
 sky130_fd_sc_hd__and2_1 _13874_ (.A(_04797_),
    .B(_04798_),
    .X(_04799_));
 sky130_fd_sc_hd__o21ba_4 _13875_ (.A1(_04678_),
    .A2(_04681_),
    .B1_N(_04679_),
    .X(_04800_));
 sky130_fd_sc_hd__a22oi_4 _13876_ (.A1(net355),
    .A2(net707),
    .B1(net716),
    .B2(net345),
    .Y(_04801_));
 sky130_fd_sc_hd__and4_1 _13877_ (.A(net345),
    .B(net355),
    .C(net708),
    .D(net716),
    .X(_04802_));
 sky130_fd_sc_hd__nor2_2 _13878_ (.A(_04801_),
    .B(_04802_),
    .Y(_04803_));
 sky130_fd_sc_hd__nand2_4 _13879_ (.A(net359),
    .B(net700),
    .Y(_04804_));
 sky130_fd_sc_hd__xnor2_4 _13880_ (.A(_04803_),
    .B(_04804_),
    .Y(_04806_));
 sky130_fd_sc_hd__and2b_1 _13881_ (.A_N(_04800_),
    .B(_04806_),
    .X(_04807_));
 sky130_fd_sc_hd__xnor2_4 _13882_ (.A(_04800_),
    .B(_04806_),
    .Y(_04808_));
 sky130_fd_sc_hd__o21ba_2 _13883_ (.A1(_04688_),
    .A2(_04691_),
    .B1_N(_04689_),
    .X(_04809_));
 sky130_fd_sc_hd__and2b_1 _13884_ (.A_N(_04809_),
    .B(_04808_),
    .X(_04810_));
 sky130_fd_sc_hd__xor2_4 _13885_ (.A(_04808_),
    .B(_04809_),
    .X(_04811_));
 sky130_fd_sc_hd__o21ba_2 _13886_ (.A1(_04694_),
    .A2(_04697_),
    .B1_N(_04693_),
    .X(_04812_));
 sky130_fd_sc_hd__nor2_4 _13887_ (.A(_04811_),
    .B(_04812_),
    .Y(_04813_));
 sky130_fd_sc_hd__and2_1 _13888_ (.A(_04811_),
    .B(_04812_),
    .X(_04814_));
 sky130_fd_sc_hd__nor2_1 _13889_ (.A(_04813_),
    .B(_04814_),
    .Y(_04815_));
 sky130_fd_sc_hd__nand2_1 _13890_ (.A(_04700_),
    .B(_04815_),
    .Y(_04817_));
 sky130_fd_sc_hd__or2_1 _13891_ (.A(_04700_),
    .B(_04815_),
    .X(_04818_));
 sky130_fd_sc_hd__nand2_1 _13892_ (.A(_04817_),
    .B(_04818_),
    .Y(_04819_));
 sky130_fd_sc_hd__nand2_8 _13893_ (.A(net377),
    .B(net681),
    .Y(_04820_));
 sky130_fd_sc_hd__a21boi_1 _13894_ (.A1(net369),
    .A2(net692),
    .B1_N(_04820_),
    .Y(_04821_));
 sky130_fd_sc_hd__and4_1 _13895_ (.A(net369),
    .B(net377),
    .C(net682),
    .D(net692),
    .X(_04822_));
 sky130_fd_sc_hd__nor2_2 _13896_ (.A(_04821_),
    .B(_04822_),
    .Y(_04823_));
 sky130_fd_sc_hd__nand2_1 _13897_ (.A(net384),
    .B(net670),
    .Y(_04824_));
 sky130_fd_sc_hd__xnor2_2 _13898_ (.A(_04823_),
    .B(_04824_),
    .Y(_04825_));
 sky130_fd_sc_hd__o21ba_1 _13899_ (.A1(_04705_),
    .A2(_04709_),
    .B1_N(_04706_),
    .X(_04826_));
 sky130_fd_sc_hd__nand2b_1 _13900_ (.A_N(_04825_),
    .B(_04826_),
    .Y(_04828_));
 sky130_fd_sc_hd__nand2b_2 _13901_ (.A_N(_04826_),
    .B(_04825_),
    .Y(_04829_));
 sky130_fd_sc_hd__nand2_2 _13902_ (.A(_04828_),
    .B(_04829_),
    .Y(_04830_));
 sky130_fd_sc_hd__nand2_2 _13903_ (.A(net392),
    .B(net662),
    .Y(_04831_));
 sky130_fd_sc_hd__xnor2_1 _13904_ (.A(_04830_),
    .B(_04831_),
    .Y(_04832_));
 sky130_fd_sc_hd__a21oi_2 _13905_ (.A1(_04712_),
    .A2(_04714_),
    .B1(_04832_),
    .Y(_04833_));
 sky130_fd_sc_hd__and3_1 _13906_ (.A(_04712_),
    .B(_04714_),
    .C(_04832_),
    .X(_04834_));
 sky130_fd_sc_hd__nor2_1 _13907_ (.A(_04833_),
    .B(_04834_),
    .Y(_04835_));
 sky130_fd_sc_hd__and3_1 _13908_ (.A(net400),
    .B(\cla_inst.in1[27] ),
    .C(_04835_),
    .X(_04836_));
 sky130_fd_sc_hd__a21oi_1 _13909_ (.A1(net400),
    .A2(net655),
    .B1(_04835_),
    .Y(_04837_));
 sky130_fd_sc_hd__or2_1 _13910_ (.A(_04836_),
    .B(_04837_),
    .X(_04839_));
 sky130_fd_sc_hd__or2_2 _13911_ (.A(_04819_),
    .B(_04839_),
    .X(_04840_));
 sky130_fd_sc_hd__nand2_1 _13912_ (.A(_04819_),
    .B(_04839_),
    .Y(_04841_));
 sky130_fd_sc_hd__and2_1 _13913_ (.A(_04840_),
    .B(_04841_),
    .X(_04842_));
 sky130_fd_sc_hd__o21a_1 _13914_ (.A1(_04703_),
    .A2(_04723_),
    .B1(_04842_),
    .X(_04843_));
 sky130_fd_sc_hd__nor3_1 _13915_ (.A(_04703_),
    .B(_04723_),
    .C(_04842_),
    .Y(_04844_));
 sky130_fd_sc_hd__nor2_1 _13916_ (.A(_04843_),
    .B(_04844_),
    .Y(_04845_));
 sky130_fd_sc_hd__nand2_1 _13917_ (.A(_04799_),
    .B(_04845_),
    .Y(_04846_));
 sky130_fd_sc_hd__or2_1 _13918_ (.A(_04799_),
    .B(_04845_),
    .X(_04847_));
 sky130_fd_sc_hd__nand2_2 _13919_ (.A(_04846_),
    .B(_04847_),
    .Y(_04848_));
 sky130_fd_sc_hd__a21o_1 _13920_ (.A1(_04684_),
    .A2(_04731_),
    .B1(_04848_),
    .X(_04850_));
 sky130_fd_sc_hd__nand3_1 _13921_ (.A(_04684_),
    .B(_04731_),
    .C(_04848_),
    .Y(_04851_));
 sky130_fd_sc_hd__nand2_2 _13922_ (.A(_04850_),
    .B(_04851_),
    .Y(_04852_));
 sky130_fd_sc_hd__xor2_2 _13923_ (.A(_04727_),
    .B(_04852_),
    .X(_04853_));
 sky130_fd_sc_hd__a21o_2 _13924_ (.A1(_04733_),
    .A2(_04736_),
    .B1(_04853_),
    .X(_04854_));
 sky130_fd_sc_hd__nand3_2 _13925_ (.A(_04733_),
    .B(_04736_),
    .C(_04853_),
    .Y(_04855_));
 sky130_fd_sc_hd__nand2_4 _13926_ (.A(_04854_),
    .B(_04855_),
    .Y(_04856_));
 sky130_fd_sc_hd__a31o_4 _13927_ (.A1(net400),
    .A2(net662),
    .A3(_04720_),
    .B1(_04717_),
    .X(_04857_));
 sky130_fd_sc_hd__nand2b_1 _13928_ (.A_N(_04856_),
    .B(_04857_),
    .Y(_04858_));
 sky130_fd_sc_hd__xor2_4 _13929_ (.A(_04856_),
    .B(_04857_),
    .X(_04859_));
 sky130_fd_sc_hd__nor2_4 _13930_ (.A(_04739_),
    .B(_04743_),
    .Y(_04861_));
 sky130_fd_sc_hd__nor2_2 _13931_ (.A(_04859_),
    .B(_04861_),
    .Y(_04862_));
 sky130_fd_sc_hd__xnor2_4 _13932_ (.A(_04859_),
    .B(_04861_),
    .Y(_04863_));
 sky130_fd_sc_hd__or2_1 _13933_ (.A(_04639_),
    .B(_04748_),
    .X(_04864_));
 sky130_fd_sc_hd__nor2_1 _13934_ (.A(_04641_),
    .B(_04864_),
    .Y(_04865_));
 sky130_fd_sc_hd__nor3b_2 _13935_ (.A(_04641_),
    .B(_04864_),
    .C_N(_04403_),
    .Y(_04866_));
 sky130_fd_sc_hd__nor3b_1 _13936_ (.A(_04639_),
    .B(_04748_),
    .C_N(_04640_),
    .Y(_04867_));
 sky130_fd_sc_hd__a211o_2 _13937_ (.A1(_04637_),
    .A2(_04746_),
    .B1(_04747_),
    .C1(_04867_),
    .X(_04868_));
 sky130_fd_sc_hd__a311oi_4 _13938_ (.A1(_03854_),
    .A2(_04404_),
    .A3(_04865_),
    .B1(_04866_),
    .C1(_04868_),
    .Y(_04869_));
 sky130_fd_sc_hd__inv_2 _13939_ (.A(net115),
    .Y(_04870_));
 sky130_fd_sc_hd__and2_1 _13940_ (.A(_04863_),
    .B(_04869_),
    .X(_04872_));
 sky130_fd_sc_hd__nor2_1 _13941_ (.A(_04863_),
    .B(_04869_),
    .Y(_04873_));
 sky130_fd_sc_hd__o31ai_1 _13942_ (.A1(net255),
    .A2(_04872_),
    .A3(_04873_),
    .B1(_04764_),
    .Y(_08659_));
 sky130_fd_sc_hd__mux2_4 _13943_ (.A0(_02639_),
    .A1(_02649_),
    .S(net552),
    .X(_04874_));
 sky130_fd_sc_hd__o21a_1 _13944_ (.A1(_02617_),
    .A2(net204),
    .B1(net205),
    .X(_04875_));
 sky130_fd_sc_hd__a21oi_4 _13945_ (.A1(net540),
    .A2(_04874_),
    .B1(_04875_),
    .Y(_04876_));
 sky130_fd_sc_hd__a22oi_2 _13946_ (.A1(net425),
    .A2(net623),
    .B1(net640),
    .B2(net409),
    .Y(_04877_));
 sky130_fd_sc_hd__nand2_2 _13947_ (.A(net408),
    .B(net623),
    .Y(_04878_));
 sky130_fd_sc_hd__and4_2 _13948_ (.A(net409),
    .B(net425),
    .C(net623),
    .D(net640),
    .X(_04879_));
 sky130_fd_sc_hd__nor2_2 _13949_ (.A(_04877_),
    .B(_04879_),
    .Y(_04880_));
 sky130_fd_sc_hd__nand2_2 _13950_ (.A(net415),
    .B(net630),
    .Y(_04882_));
 sky130_fd_sc_hd__xnor2_1 _13951_ (.A(_04880_),
    .B(_04882_),
    .Y(_04883_));
 sky130_fd_sc_hd__o21a_1 _13952_ (.A1(_04766_),
    .A2(_04769_),
    .B1(_04883_),
    .X(_04884_));
 sky130_fd_sc_hd__clkinv_2 _13953_ (.A(_04884_),
    .Y(_04885_));
 sky130_fd_sc_hd__or3_1 _13954_ (.A(_04766_),
    .B(_04769_),
    .C(_04883_),
    .X(_04886_));
 sky130_fd_sc_hd__and2_1 _13955_ (.A(_04885_),
    .B(_04886_),
    .X(_04887_));
 sky130_fd_sc_hd__nor2_1 _13956_ (.A(_04773_),
    .B(_04775_),
    .Y(_04888_));
 sky130_fd_sc_hd__o21a_1 _13957_ (.A1(_04773_),
    .A2(_04775_),
    .B1(_04887_),
    .X(_04889_));
 sky130_fd_sc_hd__nor3_1 _13958_ (.A(_04773_),
    .B(_04775_),
    .C(_04887_),
    .Y(_04890_));
 sky130_fd_sc_hd__nor2_1 _13959_ (.A(_04889_),
    .B(_04890_),
    .Y(_04891_));
 sky130_fd_sc_hd__o21ai_2 _13960_ (.A1(_04778_),
    .A2(_04780_),
    .B1(_04891_),
    .Y(_04893_));
 sky130_fd_sc_hd__or3_1 _13961_ (.A(_04778_),
    .B(_04780_),
    .C(_04891_),
    .X(_04894_));
 sky130_fd_sc_hd__and2_2 _13962_ (.A(_04893_),
    .B(_04894_),
    .X(_04895_));
 sky130_fd_sc_hd__nand2b_1 _13963_ (.A_N(_04784_),
    .B(_04895_),
    .Y(_04896_));
 sky130_fd_sc_hd__xnor2_2 _13964_ (.A(_04784_),
    .B(_04895_),
    .Y(_04897_));
 sky130_fd_sc_hd__a22oi_2 _13965_ (.A1(net331),
    .A2(net728),
    .B1(net735),
    .B2(net322),
    .Y(_04898_));
 sky130_fd_sc_hd__and4_1 _13966_ (.A(net322),
    .B(net332),
    .C(net728),
    .D(net735),
    .X(_04899_));
 sky130_fd_sc_hd__nor2_1 _13967_ (.A(_04898_),
    .B(_04899_),
    .Y(_04900_));
 sky130_fd_sc_hd__nand2_1 _13968_ (.A(net338),
    .B(net717),
    .Y(_04901_));
 sky130_fd_sc_hd__xnor2_1 _13969_ (.A(_04900_),
    .B(_04901_),
    .Y(_04902_));
 sky130_fd_sc_hd__nand2_2 _13970_ (.A(_04897_),
    .B(_04902_),
    .Y(_04904_));
 sky130_fd_sc_hd__or2_2 _13971_ (.A(_04897_),
    .B(_04902_),
    .X(_04905_));
 sky130_fd_sc_hd__nand2_4 _13972_ (.A(_04904_),
    .B(_04905_),
    .Y(_04906_));
 sky130_fd_sc_hd__a21oi_4 _13973_ (.A1(_04787_),
    .A2(_04793_),
    .B1(_04786_),
    .Y(_04907_));
 sky130_fd_sc_hd__xnor2_4 _13974_ (.A(_04906_),
    .B(_04907_),
    .Y(_04908_));
 sky130_fd_sc_hd__o21ba_4 _13975_ (.A1(_04789_),
    .A2(_04792_),
    .B1_N(_04790_),
    .X(_04909_));
 sky130_fd_sc_hd__a22oi_4 _13976_ (.A1(net355),
    .A2(net698),
    .B1(net707),
    .B2(net346),
    .Y(_04910_));
 sky130_fd_sc_hd__and4_1 _13977_ (.A(net346),
    .B(net355),
    .C(net698),
    .D(net707),
    .X(_04911_));
 sky130_fd_sc_hd__nor2_2 _13978_ (.A(_04910_),
    .B(_04911_),
    .Y(_04912_));
 sky130_fd_sc_hd__nand2_4 _13979_ (.A(net359),
    .B(net690),
    .Y(_04913_));
 sky130_fd_sc_hd__xnor2_4 _13980_ (.A(_04912_),
    .B(_04913_),
    .Y(_04915_));
 sky130_fd_sc_hd__and2b_1 _13981_ (.A_N(_04909_),
    .B(_04915_),
    .X(_04916_));
 sky130_fd_sc_hd__xnor2_4 _13982_ (.A(_04909_),
    .B(_04915_),
    .Y(_04917_));
 sky130_fd_sc_hd__o21ba_2 _13983_ (.A1(_04801_),
    .A2(_04804_),
    .B1_N(_04802_),
    .X(_04918_));
 sky130_fd_sc_hd__and2b_1 _13984_ (.A_N(_04918_),
    .B(_04917_),
    .X(_04919_));
 sky130_fd_sc_hd__xor2_4 _13985_ (.A(_04917_),
    .B(_04918_),
    .X(_04920_));
 sky130_fd_sc_hd__nor2_2 _13986_ (.A(_04807_),
    .B(_04810_),
    .Y(_04921_));
 sky130_fd_sc_hd__nor2_4 _13987_ (.A(_04920_),
    .B(_04921_),
    .Y(_04922_));
 sky130_fd_sc_hd__and2_1 _13988_ (.A(_04920_),
    .B(_04921_),
    .X(_04923_));
 sky130_fd_sc_hd__nor2_4 _13989_ (.A(_04922_),
    .B(_04923_),
    .Y(_04924_));
 sky130_fd_sc_hd__xor2_4 _13990_ (.A(_04813_),
    .B(_04924_),
    .X(_04926_));
 sky130_fd_sc_hd__a22o_1 _13991_ (.A1(net377),
    .A2(net675),
    .B1(net682),
    .B2(net369),
    .X(_04927_));
 sky130_fd_sc_hd__and2_4 _13992_ (.A(net370),
    .B(net674),
    .X(_04928_));
 sky130_fd_sc_hd__nand2_4 _13993_ (.A(net370),
    .B(net674),
    .Y(_04929_));
 sky130_fd_sc_hd__o21a_1 _13994_ (.A1(_04820_),
    .A2(_04929_),
    .B1(_04927_),
    .X(_04930_));
 sky130_fd_sc_hd__and2_1 _13995_ (.A(net385),
    .B(net663),
    .X(_04931_));
 sky130_fd_sc_hd__nor2_1 _13996_ (.A(_04930_),
    .B(_04931_),
    .Y(_04932_));
 sky130_fd_sc_hd__and2_1 _13997_ (.A(_04930_),
    .B(_04931_),
    .X(_04933_));
 sky130_fd_sc_hd__nor2_2 _13998_ (.A(_04932_),
    .B(_04933_),
    .Y(_04934_));
 sky130_fd_sc_hd__a31o_2 _13999_ (.A1(net385),
    .A2(net675),
    .A3(_04823_),
    .B1(_04822_),
    .X(_04935_));
 sky130_fd_sc_hd__nand2_1 _14000_ (.A(_04934_),
    .B(_04935_),
    .Y(_04937_));
 sky130_fd_sc_hd__xor2_2 _14001_ (.A(_04934_),
    .B(_04935_),
    .X(_04938_));
 sky130_fd_sc_hd__nand3_2 _14002_ (.A(net394),
    .B(net655),
    .C(_04938_),
    .Y(_04939_));
 sky130_fd_sc_hd__a21o_1 _14003_ (.A1(net394),
    .A2(net655),
    .B1(_04938_),
    .X(_04940_));
 sky130_fd_sc_hd__nand2_2 _14004_ (.A(_04939_),
    .B(_04940_),
    .Y(_04941_));
 sky130_fd_sc_hd__o21ai_4 _14005_ (.A1(_04830_),
    .A2(_04831_),
    .B1(_04829_),
    .Y(_04942_));
 sky130_fd_sc_hd__nand2b_1 _14006_ (.A_N(_04941_),
    .B(_04942_),
    .Y(_04943_));
 sky130_fd_sc_hd__xnor2_2 _14007_ (.A(_04941_),
    .B(_04942_),
    .Y(_04944_));
 sky130_fd_sc_hd__nand3_2 _14008_ (.A(net401),
    .B(net645),
    .C(_04944_),
    .Y(_04945_));
 sky130_fd_sc_hd__a21o_1 _14009_ (.A1(net400),
    .A2(net645),
    .B1(_04944_),
    .X(_04946_));
 sky130_fd_sc_hd__and2_1 _14010_ (.A(_04945_),
    .B(_04946_),
    .X(_04948_));
 sky130_fd_sc_hd__xnor2_2 _14011_ (.A(_04926_),
    .B(_04948_),
    .Y(_04949_));
 sky130_fd_sc_hd__a21oi_1 _14012_ (.A1(_04817_),
    .A2(_04840_),
    .B1(_04949_),
    .Y(_04950_));
 sky130_fd_sc_hd__and3_1 _14013_ (.A(_04817_),
    .B(_04840_),
    .C(_04949_),
    .X(_04951_));
 sky130_fd_sc_hd__nor2_1 _14014_ (.A(_04950_),
    .B(_04951_),
    .Y(_04952_));
 sky130_fd_sc_hd__or3_1 _14015_ (.A(_04908_),
    .B(_04950_),
    .C(_04951_),
    .X(_04953_));
 sky130_fd_sc_hd__xor2_2 _14016_ (.A(_04908_),
    .B(_04952_),
    .X(_04954_));
 sky130_fd_sc_hd__a21o_1 _14017_ (.A1(_04797_),
    .A2(_04846_),
    .B1(_04954_),
    .X(_04955_));
 sky130_fd_sc_hd__nand3_1 _14018_ (.A(_04797_),
    .B(_04846_),
    .C(_04954_),
    .Y(_04956_));
 sky130_fd_sc_hd__and2_1 _14019_ (.A(_04955_),
    .B(_04956_),
    .X(_04957_));
 sky130_fd_sc_hd__nand2_1 _14020_ (.A(_04843_),
    .B(_04957_),
    .Y(_04959_));
 sky130_fd_sc_hd__or2_1 _14021_ (.A(_04843_),
    .B(_04957_),
    .X(_04960_));
 sky130_fd_sc_hd__nand2_1 _14022_ (.A(_04959_),
    .B(_04960_),
    .Y(_04961_));
 sky130_fd_sc_hd__o31a_2 _14023_ (.A1(_04725_),
    .A2(_04726_),
    .A3(_04852_),
    .B1(_04850_),
    .X(_04962_));
 sky130_fd_sc_hd__nor2_1 _14024_ (.A(_04961_),
    .B(_04962_),
    .Y(_04963_));
 sky130_fd_sc_hd__xnor2_1 _14025_ (.A(_04961_),
    .B(_04962_),
    .Y(_04964_));
 sky130_fd_sc_hd__o21ba_1 _14026_ (.A1(_04833_),
    .A2(_04836_),
    .B1_N(_04964_),
    .X(_04965_));
 sky130_fd_sc_hd__or3b_1 _14027_ (.A(_04833_),
    .B(_04836_),
    .C_N(_04964_),
    .X(_04966_));
 sky130_fd_sc_hd__nand2b_1 _14028_ (.A_N(_04965_),
    .B(_04966_),
    .Y(_04967_));
 sky130_fd_sc_hd__a21oi_1 _14029_ (.A1(_04854_),
    .A2(_04858_),
    .B1(_04967_),
    .Y(_04968_));
 sky130_fd_sc_hd__nand3_2 _14030_ (.A(_04854_),
    .B(_04858_),
    .C(_04967_),
    .Y(_04970_));
 sky130_fd_sc_hd__nand2b_2 _14031_ (.A_N(_04968_),
    .B(_04970_),
    .Y(_04971_));
 sky130_fd_sc_hd__nor2_1 _14032_ (.A(_04862_),
    .B(_04873_),
    .Y(_04972_));
 sky130_fd_sc_hd__or2_1 _14033_ (.A(_04971_),
    .B(_04972_),
    .X(_04973_));
 sky130_fd_sc_hd__nand2_1 _14034_ (.A(_04971_),
    .B(_04972_),
    .Y(_04974_));
 sky130_fd_sc_hd__a31o_1 _14035_ (.A1(net258),
    .A2(_04973_),
    .A3(_04974_),
    .B1(_04876_),
    .X(_08660_));
 sky130_fd_sc_hd__mux2_4 _14036_ (.A0(_02851_),
    .A1(_02857_),
    .S(net552),
    .X(_04975_));
 sky130_fd_sc_hd__o21a_1 _14037_ (.A1(_02832_),
    .A2(net204),
    .B1(net205),
    .X(_04976_));
 sky130_fd_sc_hd__a21oi_4 _14038_ (.A1(net540),
    .A2(_04975_),
    .B1(_04976_),
    .Y(_04977_));
 sky130_fd_sc_hd__a31o_4 _14039_ (.A1(net415),
    .A2(net631),
    .A3(_04880_),
    .B1(_04879_),
    .X(_04978_));
 sky130_fd_sc_hd__a22o_1 _14040_ (.A1(net416),
    .A2(net623),
    .B1(net631),
    .B2(net408),
    .X(_04980_));
 sky130_fd_sc_hd__o21a_2 _14041_ (.A1(_04878_),
    .A2(_04882_),
    .B1(_04980_),
    .X(_04981_));
 sky130_fd_sc_hd__nand2_2 _14042_ (.A(_04978_),
    .B(_04981_),
    .Y(_04982_));
 sky130_fd_sc_hd__xnor2_4 _14043_ (.A(_04978_),
    .B(_04981_),
    .Y(_04983_));
 sky130_fd_sc_hd__nor2_1 _14044_ (.A(_04884_),
    .B(_04889_),
    .Y(_04984_));
 sky130_fd_sc_hd__xnor2_1 _14045_ (.A(_04983_),
    .B(_04984_),
    .Y(_04985_));
 sky130_fd_sc_hd__nor2_1 _14046_ (.A(_04893_),
    .B(_04985_),
    .Y(_04986_));
 sky130_fd_sc_hd__and2_1 _14047_ (.A(_04893_),
    .B(_04985_),
    .X(_04987_));
 sky130_fd_sc_hd__or2_4 _14048_ (.A(_04986_),
    .B(_04987_),
    .X(_04988_));
 sky130_fd_sc_hd__a22oi_1 _14049_ (.A1(net331),
    .A2(net717),
    .B1(net727),
    .B2(net322),
    .Y(_04989_));
 sky130_fd_sc_hd__and4_1 _14050_ (.A(net322),
    .B(net331),
    .C(net717),
    .D(net728),
    .X(_04991_));
 sky130_fd_sc_hd__or2_1 _14051_ (.A(_04989_),
    .B(_04991_),
    .X(_04992_));
 sky130_fd_sc_hd__nand2_1 _14052_ (.A(net338),
    .B(net709),
    .Y(_04993_));
 sky130_fd_sc_hd__nor2_2 _14053_ (.A(_04992_),
    .B(_04993_),
    .Y(_04994_));
 sky130_fd_sc_hd__and2_1 _14054_ (.A(_04992_),
    .B(_04993_),
    .X(_04995_));
 sky130_fd_sc_hd__nor2_2 _14055_ (.A(_04994_),
    .B(_04995_),
    .Y(_04996_));
 sky130_fd_sc_hd__and2b_1 _14056_ (.A_N(_04988_),
    .B(_04996_),
    .X(_04997_));
 sky130_fd_sc_hd__xor2_4 _14057_ (.A(_04988_),
    .B(_04996_),
    .X(_04998_));
 sky130_fd_sc_hd__nand2_1 _14058_ (.A(_04896_),
    .B(_04904_),
    .Y(_04999_));
 sky130_fd_sc_hd__a21o_1 _14059_ (.A1(_04896_),
    .A2(_04904_),
    .B1(_04998_),
    .X(_05000_));
 sky130_fd_sc_hd__xnor2_2 _14060_ (.A(_04998_),
    .B(_04999_),
    .Y(_05002_));
 sky130_fd_sc_hd__o21ba_2 _14061_ (.A1(_04898_),
    .A2(_04901_),
    .B1_N(_04899_),
    .X(_05003_));
 sky130_fd_sc_hd__a22oi_4 _14062_ (.A1(net353),
    .A2(net691),
    .B1(net700),
    .B2(net347),
    .Y(_05004_));
 sky130_fd_sc_hd__and4_1 _14063_ (.A(net347),
    .B(net353),
    .C(net691),
    .D(net700),
    .X(_05005_));
 sky130_fd_sc_hd__nor2_1 _14064_ (.A(_05004_),
    .B(_05005_),
    .Y(_05006_));
 sky130_fd_sc_hd__nand2_2 _14065_ (.A(net360),
    .B(net682),
    .Y(_05007_));
 sky130_fd_sc_hd__xnor2_2 _14066_ (.A(_05006_),
    .B(_05007_),
    .Y(_05008_));
 sky130_fd_sc_hd__and2b_1 _14067_ (.A_N(_05003_),
    .B(_05008_),
    .X(_05009_));
 sky130_fd_sc_hd__xnor2_2 _14068_ (.A(_05003_),
    .B(_05008_),
    .Y(_05010_));
 sky130_fd_sc_hd__o21ba_2 _14069_ (.A1(_04910_),
    .A2(_04913_),
    .B1_N(_04911_),
    .X(_05011_));
 sky130_fd_sc_hd__and2b_1 _14070_ (.A_N(_05011_),
    .B(_05010_),
    .X(_05013_));
 sky130_fd_sc_hd__xor2_1 _14071_ (.A(_05010_),
    .B(_05011_),
    .X(_05014_));
 sky130_fd_sc_hd__nor2_1 _14072_ (.A(_04916_),
    .B(_04919_),
    .Y(_05015_));
 sky130_fd_sc_hd__or2_2 _14073_ (.A(_05014_),
    .B(_05015_),
    .X(_05016_));
 sky130_fd_sc_hd__nand2_1 _14074_ (.A(_05014_),
    .B(_05015_),
    .Y(_05017_));
 sky130_fd_sc_hd__and2_1 _14075_ (.A(_05016_),
    .B(_05017_),
    .X(_05018_));
 sky130_fd_sc_hd__nand2_2 _14076_ (.A(_04922_),
    .B(_05018_),
    .Y(_05019_));
 sky130_fd_sc_hd__or2_1 _14077_ (.A(_04922_),
    .B(_05018_),
    .X(_05020_));
 sky130_fd_sc_hd__nand2_1 _14078_ (.A(_05019_),
    .B(_05020_),
    .Y(_05021_));
 sky130_fd_sc_hd__a21oi_2 _14079_ (.A1(net377),
    .A2(net665),
    .B1(_04928_),
    .Y(_05022_));
 sky130_fd_sc_hd__and3_4 _14080_ (.A(net377),
    .B(net665),
    .C(_04928_),
    .X(_05024_));
 sky130_fd_sc_hd__nor2_4 _14081_ (.A(_05022_),
    .B(_05024_),
    .Y(_05025_));
 sky130_fd_sc_hd__nand2_2 _14082_ (.A(net385),
    .B(net657),
    .Y(_05026_));
 sky130_fd_sc_hd__and3_2 _14083_ (.A(net385),
    .B(net657),
    .C(_05025_),
    .X(_05027_));
 sky130_fd_sc_hd__xnor2_4 _14084_ (.A(_05025_),
    .B(_05026_),
    .Y(_05028_));
 sky130_fd_sc_hd__o21ba_1 _14085_ (.A1(_04820_),
    .A2(_04929_),
    .B1_N(_04933_),
    .X(_05029_));
 sky130_fd_sc_hd__nand2b_1 _14086_ (.A_N(_05028_),
    .B(_05029_),
    .Y(_05030_));
 sky130_fd_sc_hd__nand2b_4 _14087_ (.A_N(_05029_),
    .B(_05028_),
    .Y(_05031_));
 sky130_fd_sc_hd__nand2_4 _14088_ (.A(_05030_),
    .B(_05031_),
    .Y(_05032_));
 sky130_fd_sc_hd__nand2_2 _14089_ (.A(net394),
    .B(net645),
    .Y(_05033_));
 sky130_fd_sc_hd__xnor2_2 _14090_ (.A(_05032_),
    .B(_05033_),
    .Y(_05035_));
 sky130_fd_sc_hd__a21oi_2 _14091_ (.A1(_04937_),
    .A2(_04939_),
    .B1(_05035_),
    .Y(_05036_));
 sky130_fd_sc_hd__and3_1 _14092_ (.A(_04937_),
    .B(_04939_),
    .C(_05035_),
    .X(_05037_));
 sky130_fd_sc_hd__nor2_1 _14093_ (.A(_05036_),
    .B(_05037_),
    .Y(_05038_));
 sky130_fd_sc_hd__and3_1 _14094_ (.A(net402),
    .B(net635),
    .C(_05038_),
    .X(_05039_));
 sky130_fd_sc_hd__a21oi_1 _14095_ (.A1(net402),
    .A2(net635),
    .B1(_05038_),
    .Y(_05040_));
 sky130_fd_sc_hd__or2_1 _14096_ (.A(_05039_),
    .B(_05040_),
    .X(_05041_));
 sky130_fd_sc_hd__or2_4 _14097_ (.A(_05021_),
    .B(_05041_),
    .X(_05042_));
 sky130_fd_sc_hd__nand2_1 _14098_ (.A(_05021_),
    .B(_05041_),
    .Y(_05043_));
 sky130_fd_sc_hd__nand2_1 _14099_ (.A(_05042_),
    .B(_05043_),
    .Y(_05044_));
 sky130_fd_sc_hd__a32o_2 _14100_ (.A1(_04926_),
    .A2(_04945_),
    .A3(_04946_),
    .B1(_04924_),
    .B2(_04813_),
    .X(_05046_));
 sky130_fd_sc_hd__and3_1 _14101_ (.A(_05042_),
    .B(_05043_),
    .C(_05046_),
    .X(_05047_));
 sky130_fd_sc_hd__xnor2_1 _14102_ (.A(_05044_),
    .B(_05046_),
    .Y(_05048_));
 sky130_fd_sc_hd__nand2_1 _14103_ (.A(_05002_),
    .B(_05048_),
    .Y(_05049_));
 sky130_fd_sc_hd__or2_1 _14104_ (.A(_05002_),
    .B(_05048_),
    .X(_05050_));
 sky130_fd_sc_hd__nand2_2 _14105_ (.A(_05049_),
    .B(_05050_),
    .Y(_05051_));
 sky130_fd_sc_hd__o21ai_2 _14106_ (.A1(_04906_),
    .A2(_04907_),
    .B1(_04953_),
    .Y(_05052_));
 sky130_fd_sc_hd__nand2b_1 _14107_ (.A_N(_05051_),
    .B(_05052_),
    .Y(_05053_));
 sky130_fd_sc_hd__xor2_2 _14108_ (.A(_05051_),
    .B(_05052_),
    .X(_05054_));
 sky130_fd_sc_hd__a211o_2 _14109_ (.A1(_04817_),
    .A2(_04840_),
    .B1(_04949_),
    .C1(_05054_),
    .X(_05055_));
 sky130_fd_sc_hd__nand2b_1 _14110_ (.A_N(_04950_),
    .B(_05054_),
    .Y(_05057_));
 sky130_fd_sc_hd__nand2_1 _14111_ (.A(_05055_),
    .B(_05057_),
    .Y(_05058_));
 sky130_fd_sc_hd__a21o_1 _14112_ (.A1(_04955_),
    .A2(_04959_),
    .B1(_05058_),
    .X(_05059_));
 sky130_fd_sc_hd__nand3_1 _14113_ (.A(_04955_),
    .B(_04959_),
    .C(_05058_),
    .Y(_05060_));
 sky130_fd_sc_hd__nand2_1 _14114_ (.A(_05059_),
    .B(_05060_),
    .Y(_05061_));
 sky130_fd_sc_hd__nand2_1 _14115_ (.A(_04943_),
    .B(_04945_),
    .Y(_05062_));
 sky130_fd_sc_hd__nand2b_1 _14116_ (.A_N(_05061_),
    .B(_05062_),
    .Y(_05063_));
 sky130_fd_sc_hd__xor2_1 _14117_ (.A(_05061_),
    .B(_05062_),
    .X(_05064_));
 sky130_fd_sc_hd__o21ba_1 _14118_ (.A1(_04963_),
    .A2(_04965_),
    .B1_N(_05064_),
    .X(_05065_));
 sky130_fd_sc_hd__or3b_1 _14119_ (.A(_04963_),
    .B(_04965_),
    .C_N(_05064_),
    .X(_05066_));
 sky130_fd_sc_hd__nand2b_1 _14120_ (.A_N(_05065_),
    .B(_05066_),
    .Y(_05068_));
 sky130_fd_sc_hd__o21a_1 _14121_ (.A1(_04862_),
    .A2(_04968_),
    .B1(_04970_),
    .X(_05069_));
 sky130_fd_sc_hd__nor2_1 _14122_ (.A(_04863_),
    .B(_04971_),
    .Y(_05070_));
 sky130_fd_sc_hd__a21oi_1 _14123_ (.A1(_04870_),
    .A2(_05070_),
    .B1(_05069_),
    .Y(_05071_));
 sky130_fd_sc_hd__nand2_1 _14124_ (.A(_05068_),
    .B(_05071_),
    .Y(_05072_));
 sky130_fd_sc_hd__or2_1 _14125_ (.A(_05068_),
    .B(_05071_),
    .X(_05073_));
 sky130_fd_sc_hd__a31o_1 _14126_ (.A1(net258),
    .A2(_05072_),
    .A3(_05073_),
    .B1(_04977_),
    .X(_08661_));
 sky130_fd_sc_hd__mux2_4 _14127_ (.A0(_03019_),
    .A1(_03022_),
    .S(net554),
    .X(_05074_));
 sky130_fd_sc_hd__o21a_1 _14128_ (.A1(_03012_),
    .A2(net204),
    .B1(net205),
    .X(_05075_));
 sky130_fd_sc_hd__a21oi_4 _14129_ (.A1(net540),
    .A2(_05074_),
    .B1(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hd__nor3b_1 _14130_ (.A(_04888_),
    .B(_04983_),
    .C_N(_04887_),
    .Y(_05078_));
 sky130_fd_sc_hd__inv_2 _14131_ (.A(_05078_),
    .Y(_05079_));
 sky130_fd_sc_hd__a21oi_4 _14132_ (.A1(_04882_),
    .A2(_04982_),
    .B1(_04878_),
    .Y(_05080_));
 sky130_fd_sc_hd__a21o_1 _14133_ (.A1(_04878_),
    .A2(_04982_),
    .B1(_05080_),
    .X(_05081_));
 sky130_fd_sc_hd__nor3_4 _14134_ (.A(_04885_),
    .B(_04983_),
    .C(_05081_),
    .Y(_05082_));
 sky130_fd_sc_hd__o21a_1 _14135_ (.A1(_04885_),
    .A2(_04983_),
    .B1(_05081_),
    .X(_05083_));
 sky130_fd_sc_hd__or2_1 _14136_ (.A(_05082_),
    .B(_05083_),
    .X(_05084_));
 sky130_fd_sc_hd__nor2_2 _14137_ (.A(_05079_),
    .B(_05084_),
    .Y(_05085_));
 sky130_fd_sc_hd__and2_1 _14138_ (.A(_05079_),
    .B(_05084_),
    .X(_05086_));
 sky130_fd_sc_hd__or2_1 _14139_ (.A(_05085_),
    .B(_05086_),
    .X(_05087_));
 sky130_fd_sc_hd__a22oi_1 _14140_ (.A1(net331),
    .A2(net709),
    .B1(net717),
    .B2(net321),
    .Y(_05089_));
 sky130_fd_sc_hd__and4_1 _14141_ (.A(net322),
    .B(net331),
    .C(net709),
    .D(net717),
    .X(_05090_));
 sky130_fd_sc_hd__or2_1 _14142_ (.A(_05089_),
    .B(_05090_),
    .X(_05091_));
 sky130_fd_sc_hd__nand2_1 _14143_ (.A(net339),
    .B(net700),
    .Y(_05092_));
 sky130_fd_sc_hd__nor2_1 _14144_ (.A(_05091_),
    .B(_05092_),
    .Y(_05093_));
 sky130_fd_sc_hd__and2_1 _14145_ (.A(_05091_),
    .B(_05092_),
    .X(_05094_));
 sky130_fd_sc_hd__nor2_1 _14146_ (.A(_05093_),
    .B(_05094_),
    .Y(_05095_));
 sky130_fd_sc_hd__and2b_1 _14147_ (.A_N(_05087_),
    .B(_05095_),
    .X(_05096_));
 sky130_fd_sc_hd__xnor2_1 _14148_ (.A(_05087_),
    .B(_05095_),
    .Y(_05097_));
 sky130_fd_sc_hd__o21a_2 _14149_ (.A1(_04986_),
    .A2(_04997_),
    .B1(_05097_),
    .X(_05098_));
 sky130_fd_sc_hd__nor3_1 _14150_ (.A(_04986_),
    .B(_04997_),
    .C(_05097_),
    .Y(_05100_));
 sky130_fd_sc_hd__nor2_2 _14151_ (.A(_05098_),
    .B(_05100_),
    .Y(_05101_));
 sky130_fd_sc_hd__a22oi_2 _14152_ (.A1(net353),
    .A2(net681),
    .B1(net691),
    .B2(net346),
    .Y(_05102_));
 sky130_fd_sc_hd__and4_1 _14153_ (.A(net346),
    .B(net353),
    .C(net681),
    .D(net692),
    .X(_05103_));
 sky130_fd_sc_hd__nor2_1 _14154_ (.A(_05102_),
    .B(_05103_),
    .Y(_05104_));
 sky130_fd_sc_hd__nand2_2 _14155_ (.A(net361),
    .B(net673),
    .Y(_05105_));
 sky130_fd_sc_hd__xnor2_2 _14156_ (.A(_05104_),
    .B(_05105_),
    .Y(_05106_));
 sky130_fd_sc_hd__o21a_1 _14157_ (.A1(_04991_),
    .A2(_04994_),
    .B1(_05106_),
    .X(_05107_));
 sky130_fd_sc_hd__nor3_2 _14158_ (.A(_04991_),
    .B(_04994_),
    .C(_05106_),
    .Y(_05108_));
 sky130_fd_sc_hd__nor2_2 _14159_ (.A(_05107_),
    .B(_05108_),
    .Y(_05109_));
 sky130_fd_sc_hd__o21ba_4 _14160_ (.A1(_05004_),
    .A2(_05007_),
    .B1_N(_05005_),
    .X(_05111_));
 sky130_fd_sc_hd__xor2_4 _14161_ (.A(_05109_),
    .B(_05111_),
    .X(_05112_));
 sky130_fd_sc_hd__nor2_4 _14162_ (.A(_05009_),
    .B(_05013_),
    .Y(_05113_));
 sky130_fd_sc_hd__xor2_2 _14163_ (.A(_05112_),
    .B(_05113_),
    .X(_05114_));
 sky130_fd_sc_hd__and2b_1 _14164_ (.A_N(_05016_),
    .B(_05114_),
    .X(_05115_));
 sky130_fd_sc_hd__xnor2_1 _14165_ (.A(_05016_),
    .B(_05114_),
    .Y(_05116_));
 sky130_fd_sc_hd__a22oi_4 _14166_ (.A1(net378),
    .A2(net657),
    .B1(net665),
    .B2(net368),
    .Y(_05117_));
 sky130_fd_sc_hd__and4_4 _14167_ (.A(net368),
    .B(net377),
    .C(net657),
    .D(net665),
    .X(_05118_));
 sky130_fd_sc_hd__nand2_2 _14168_ (.A(net385),
    .B(net650),
    .Y(_05119_));
 sky130_fd_sc_hd__o21a_1 _14169_ (.A1(_05117_),
    .A2(_05118_),
    .B1(_05119_),
    .X(_05120_));
 sky130_fd_sc_hd__nor3_4 _14170_ (.A(_05117_),
    .B(_05118_),
    .C(_05119_),
    .Y(_05122_));
 sky130_fd_sc_hd__nor2_2 _14171_ (.A(_05120_),
    .B(_05122_),
    .Y(_05123_));
 sky130_fd_sc_hd__o21ai_4 _14172_ (.A1(_05024_),
    .A2(_05027_),
    .B1(_05123_),
    .Y(_05124_));
 sky130_fd_sc_hd__or3_1 _14173_ (.A(_05024_),
    .B(_05027_),
    .C(_05123_),
    .X(_05125_));
 sky130_fd_sc_hd__and2_4 _14174_ (.A(_05124_),
    .B(_05125_),
    .X(_05126_));
 sky130_fd_sc_hd__nand2_2 _14175_ (.A(net394),
    .B(net640),
    .Y(_05127_));
 sky130_fd_sc_hd__nand3_2 _14176_ (.A(net394),
    .B(net640),
    .C(_05126_),
    .Y(_05128_));
 sky130_fd_sc_hd__xor2_4 _14177_ (.A(_05126_),
    .B(_05127_),
    .X(_05129_));
 sky130_fd_sc_hd__o21ai_4 _14178_ (.A1(_05032_),
    .A2(_05033_),
    .B1(_05031_),
    .Y(_05130_));
 sky130_fd_sc_hd__nand2b_1 _14179_ (.A_N(_05129_),
    .B(_05130_),
    .Y(_05131_));
 sky130_fd_sc_hd__xnor2_2 _14180_ (.A(_05129_),
    .B(_05130_),
    .Y(_05133_));
 sky130_fd_sc_hd__nand3_2 _14181_ (.A(net402),
    .B(net631),
    .C(_05133_),
    .Y(_05134_));
 sky130_fd_sc_hd__a21o_1 _14182_ (.A1(\cla_inst.in2[21] ),
    .A2(net631),
    .B1(_05133_),
    .X(_05135_));
 sky130_fd_sc_hd__and2_1 _14183_ (.A(_05134_),
    .B(_05135_),
    .X(_05136_));
 sky130_fd_sc_hd__and3_1 _14184_ (.A(_05116_),
    .B(_05134_),
    .C(_05135_),
    .X(_05137_));
 sky130_fd_sc_hd__nor2_1 _14185_ (.A(_05116_),
    .B(_05136_),
    .Y(_05138_));
 sky130_fd_sc_hd__or2_2 _14186_ (.A(_05137_),
    .B(_05138_),
    .X(_05139_));
 sky130_fd_sc_hd__a21oi_4 _14187_ (.A1(_05019_),
    .A2(_05042_),
    .B1(_05139_),
    .Y(_05140_));
 sky130_fd_sc_hd__and3_1 _14188_ (.A(_05019_),
    .B(_05042_),
    .C(_05139_),
    .X(_05141_));
 sky130_fd_sc_hd__nor2_2 _14189_ (.A(_05140_),
    .B(_05141_),
    .Y(_05142_));
 sky130_fd_sc_hd__xnor2_2 _14190_ (.A(_05101_),
    .B(_05142_),
    .Y(_05144_));
 sky130_fd_sc_hd__a21o_1 _14191_ (.A1(_05000_),
    .A2(_05049_),
    .B1(_05144_),
    .X(_05145_));
 sky130_fd_sc_hd__nand3_1 _14192_ (.A(_05000_),
    .B(_05049_),
    .C(_05144_),
    .Y(_05146_));
 sky130_fd_sc_hd__nand2_2 _14193_ (.A(_05145_),
    .B(_05146_),
    .Y(_05147_));
 sky130_fd_sc_hd__or3b_2 _14194_ (.A(_05044_),
    .B(_05147_),
    .C_N(_05046_),
    .X(_05148_));
 sky130_fd_sc_hd__xor2_2 _14195_ (.A(_05047_),
    .B(_05147_),
    .X(_05149_));
 sky130_fd_sc_hd__a21oi_2 _14196_ (.A1(_05053_),
    .A2(_05055_),
    .B1(_05149_),
    .Y(_05150_));
 sky130_fd_sc_hd__and3_1 _14197_ (.A(_05053_),
    .B(_05055_),
    .C(_05149_),
    .X(_05151_));
 sky130_fd_sc_hd__or2_1 _14198_ (.A(_05150_),
    .B(_05151_),
    .X(_05152_));
 sky130_fd_sc_hd__o21ba_1 _14199_ (.A1(_05036_),
    .A2(_05039_),
    .B1_N(_05152_),
    .X(_05153_));
 sky130_fd_sc_hd__or3b_1 _14200_ (.A(_05036_),
    .B(_05039_),
    .C_N(_05152_),
    .X(_05155_));
 sky130_fd_sc_hd__nand2b_1 _14201_ (.A_N(_05153_),
    .B(_05155_),
    .Y(_05156_));
 sky130_fd_sc_hd__and3_1 _14202_ (.A(_05059_),
    .B(_05063_),
    .C(_05156_),
    .X(_05157_));
 sky130_fd_sc_hd__a21oi_1 _14203_ (.A1(_05059_),
    .A2(_05063_),
    .B1(_05156_),
    .Y(_05158_));
 sky130_fd_sc_hd__or2_1 _14204_ (.A(_05157_),
    .B(_05158_),
    .X(_05159_));
 sky130_fd_sc_hd__and2b_1 _14205_ (.A_N(_05065_),
    .B(_05073_),
    .X(_05160_));
 sky130_fd_sc_hd__nand2_1 _14206_ (.A(_05159_),
    .B(_05160_),
    .Y(_05161_));
 sky130_fd_sc_hd__or2_1 _14207_ (.A(_05159_),
    .B(_05160_),
    .X(_05162_));
 sky130_fd_sc_hd__a31o_1 _14208_ (.A1(net258),
    .A2(_05161_),
    .A3(_05162_),
    .B1(_05076_),
    .X(_08662_));
 sky130_fd_sc_hd__mux2_2 _14209_ (.A0(_03180_),
    .A1(_03194_),
    .S(net553),
    .X(_05163_));
 sky130_fd_sc_hd__or2_1 _14210_ (.A(_03188_),
    .B(net204),
    .X(_05165_));
 sky130_fd_sc_hd__a22o_2 _14211_ (.A1(net537),
    .A2(_05163_),
    .B1(_05165_),
    .B2(_03686_),
    .X(_05166_));
 sky130_fd_sc_hd__a22oi_2 _14212_ (.A1(net331),
    .A2(net700),
    .B1(net709),
    .B2(net321),
    .Y(_05167_));
 sky130_fd_sc_hd__and4_1 _14213_ (.A(net322),
    .B(net331),
    .C(net700),
    .D(net709),
    .X(_05168_));
 sky130_fd_sc_hd__nor2_1 _14214_ (.A(_05167_),
    .B(_05168_),
    .Y(_05169_));
 sky130_fd_sc_hd__nand2_2 _14215_ (.A(net339),
    .B(net692),
    .Y(_05170_));
 sky130_fd_sc_hd__xnor2_2 _14216_ (.A(_05169_),
    .B(_05170_),
    .Y(_05171_));
 sky130_fd_sc_hd__o21ai_4 _14217_ (.A1(_05080_),
    .A2(_05082_),
    .B1(_05171_),
    .Y(_05172_));
 sky130_fd_sc_hd__or3_1 _14218_ (.A(_05080_),
    .B(_05082_),
    .C(_05171_),
    .X(_05173_));
 sky130_fd_sc_hd__and2_1 _14219_ (.A(_05172_),
    .B(_05173_),
    .X(_05174_));
 sky130_fd_sc_hd__o21ai_4 _14220_ (.A1(_05085_),
    .A2(_05096_),
    .B1(_05174_),
    .Y(_05176_));
 sky130_fd_sc_hd__or3_1 _14221_ (.A(_05085_),
    .B(_05096_),
    .C(_05174_),
    .X(_05177_));
 sky130_fd_sc_hd__nand2_1 _14222_ (.A(_05176_),
    .B(_05177_),
    .Y(_05178_));
 sky130_fd_sc_hd__a22oi_2 _14223_ (.A1(net353),
    .A2(net673),
    .B1(net682),
    .B2(net347),
    .Y(_05179_));
 sky130_fd_sc_hd__and4_1 _14224_ (.A(net346),
    .B(net354),
    .C(net673),
    .D(net682),
    .X(_05180_));
 sky130_fd_sc_hd__nor2_1 _14225_ (.A(_05179_),
    .B(_05180_),
    .Y(_05181_));
 sky130_fd_sc_hd__nand2_4 _14226_ (.A(net360),
    .B(net665),
    .Y(_05182_));
 sky130_fd_sc_hd__xnor2_1 _14227_ (.A(_05181_),
    .B(_05182_),
    .Y(_05183_));
 sky130_fd_sc_hd__o21a_1 _14228_ (.A1(_05090_),
    .A2(_05093_),
    .B1(_05183_),
    .X(_05184_));
 sky130_fd_sc_hd__nor3_1 _14229_ (.A(_05090_),
    .B(_05093_),
    .C(_05183_),
    .Y(_05185_));
 sky130_fd_sc_hd__nor2_1 _14230_ (.A(_05184_),
    .B(_05185_),
    .Y(_05187_));
 sky130_fd_sc_hd__o21ba_1 _14231_ (.A1(_05102_),
    .A2(_05105_),
    .B1_N(_05103_),
    .X(_05188_));
 sky130_fd_sc_hd__xor2_1 _14232_ (.A(_05187_),
    .B(_05188_),
    .X(_05189_));
 sky130_fd_sc_hd__o21ba_1 _14233_ (.A1(_05108_),
    .A2(_05111_),
    .B1_N(_05107_),
    .X(_05190_));
 sky130_fd_sc_hd__or2_1 _14234_ (.A(_05189_),
    .B(_05190_),
    .X(_05191_));
 sky130_fd_sc_hd__nand2_1 _14235_ (.A(_05189_),
    .B(_05190_),
    .Y(_05192_));
 sky130_fd_sc_hd__and2_1 _14236_ (.A(_05191_),
    .B(_05192_),
    .X(_05193_));
 sky130_fd_sc_hd__nor3b_4 _14237_ (.A(_05112_),
    .B(_05113_),
    .C_N(_05193_),
    .Y(_05194_));
 sky130_fd_sc_hd__o21ba_1 _14238_ (.A1(_05112_),
    .A2(_05113_),
    .B1_N(_05193_),
    .X(_05195_));
 sky130_fd_sc_hd__nor2_1 _14239_ (.A(_05194_),
    .B(_05195_),
    .Y(_05196_));
 sky130_fd_sc_hd__a22oi_2 _14240_ (.A1(net377),
    .A2(net650),
    .B1(net657),
    .B2(net368),
    .Y(_05198_));
 sky130_fd_sc_hd__and4_1 _14241_ (.A(net368),
    .B(net378),
    .C(net650),
    .D(net657),
    .X(_05199_));
 sky130_fd_sc_hd__nor2_1 _14242_ (.A(_05198_),
    .B(_05199_),
    .Y(_05200_));
 sky130_fd_sc_hd__nand2_2 _14243_ (.A(net385),
    .B(net640),
    .Y(_05201_));
 sky130_fd_sc_hd__xnor2_2 _14244_ (.A(_05200_),
    .B(_05201_),
    .Y(_05202_));
 sky130_fd_sc_hd__or3_1 _14245_ (.A(_05118_),
    .B(_05122_),
    .C(_05202_),
    .X(_05203_));
 sky130_fd_sc_hd__o21ai_4 _14246_ (.A1(_05118_),
    .A2(_05122_),
    .B1(_05202_),
    .Y(_05204_));
 sky130_fd_sc_hd__and2_2 _14247_ (.A(_05203_),
    .B(_05204_),
    .X(_05205_));
 sky130_fd_sc_hd__nand3_4 _14248_ (.A(net394),
    .B(net631),
    .C(_05205_),
    .Y(_05206_));
 sky130_fd_sc_hd__a21o_1 _14249_ (.A1(net394),
    .A2(net631),
    .B1(_05205_),
    .X(_05207_));
 sky130_fd_sc_hd__nand2_2 _14250_ (.A(_05206_),
    .B(_05207_),
    .Y(_05209_));
 sky130_fd_sc_hd__a21oi_4 _14251_ (.A1(_05124_),
    .A2(_05128_),
    .B1(_05209_),
    .Y(_05210_));
 sky130_fd_sc_hd__and3_1 _14252_ (.A(_05124_),
    .B(_05128_),
    .C(_05209_),
    .X(_05211_));
 sky130_fd_sc_hd__nor2_4 _14253_ (.A(_05210_),
    .B(_05211_),
    .Y(_05212_));
 sky130_fd_sc_hd__nand2_1 _14254_ (.A(net402),
    .B(net622),
    .Y(_05213_));
 sky130_fd_sc_hd__xnor2_2 _14255_ (.A(_05212_),
    .B(_05213_),
    .Y(_05214_));
 sky130_fd_sc_hd__and2_2 _14256_ (.A(_05196_),
    .B(_05214_),
    .X(_05215_));
 sky130_fd_sc_hd__nand2_1 _14257_ (.A(_05196_),
    .B(_05214_),
    .Y(_05216_));
 sky130_fd_sc_hd__or2_1 _14258_ (.A(_05196_),
    .B(_05214_),
    .X(_05217_));
 sky130_fd_sc_hd__o211a_2 _14259_ (.A1(_05115_),
    .A2(_05137_),
    .B1(_05216_),
    .C1(_05217_),
    .X(_05218_));
 sky130_fd_sc_hd__a211oi_2 _14260_ (.A1(_05216_),
    .A2(_05217_),
    .B1(_05115_),
    .C1(_05137_),
    .Y(_05220_));
 sky130_fd_sc_hd__o21ai_1 _14261_ (.A1(_05218_),
    .A2(_05220_),
    .B1(_05178_),
    .Y(_05221_));
 sky130_fd_sc_hd__or3_4 _14262_ (.A(_05178_),
    .B(_05218_),
    .C(_05220_),
    .X(_05222_));
 sky130_fd_sc_hd__nand2_1 _14263_ (.A(_05221_),
    .B(_05222_),
    .Y(_05223_));
 sky130_fd_sc_hd__a21o_1 _14264_ (.A1(_05101_),
    .A2(_05142_),
    .B1(_05098_),
    .X(_05224_));
 sky130_fd_sc_hd__and3_1 _14265_ (.A(_05221_),
    .B(_05222_),
    .C(_05224_),
    .X(_05225_));
 sky130_fd_sc_hd__xnor2_2 _14266_ (.A(_05223_),
    .B(_05224_),
    .Y(_05226_));
 sky130_fd_sc_hd__and2_1 _14267_ (.A(_05140_),
    .B(_05226_),
    .X(_05227_));
 sky130_fd_sc_hd__xnor2_2 _14268_ (.A(_05140_),
    .B(_05226_),
    .Y(_05228_));
 sky130_fd_sc_hd__a21oi_2 _14269_ (.A1(_05145_),
    .A2(_05148_),
    .B1(_05228_),
    .Y(_05229_));
 sky130_fd_sc_hd__and3_1 _14270_ (.A(_05145_),
    .B(_05148_),
    .C(_05228_),
    .X(_05231_));
 sky130_fd_sc_hd__or2_1 _14271_ (.A(_05229_),
    .B(_05231_),
    .X(_05232_));
 sky130_fd_sc_hd__a21oi_1 _14272_ (.A1(_05131_),
    .A2(_05134_),
    .B1(_05232_),
    .Y(_05233_));
 sky130_fd_sc_hd__and3_1 _14273_ (.A(_05131_),
    .B(_05134_),
    .C(_05232_),
    .X(_05234_));
 sky130_fd_sc_hd__or2_1 _14274_ (.A(_05233_),
    .B(_05234_),
    .X(_05235_));
 sky130_fd_sc_hd__o21ba_1 _14275_ (.A1(_05150_),
    .A2(_05153_),
    .B1_N(_05235_),
    .X(_05236_));
 sky130_fd_sc_hd__or3b_1 _14276_ (.A(_05150_),
    .B(_05153_),
    .C_N(_05235_),
    .X(_05237_));
 sky130_fd_sc_hd__nand2b_1 _14277_ (.A_N(_05236_),
    .B(_05237_),
    .Y(_05238_));
 sky130_fd_sc_hd__nor2_1 _14278_ (.A(_05068_),
    .B(_05159_),
    .Y(_05239_));
 sky130_fd_sc_hd__nor2_1 _14279_ (.A(_05065_),
    .B(_05158_),
    .Y(_05240_));
 sky130_fd_sc_hd__o2bb2a_1 _14280_ (.A1_N(_05069_),
    .A2_N(_05239_),
    .B1(_05240_),
    .B2(_05157_),
    .X(_05242_));
 sky130_fd_sc_hd__nand2_2 _14281_ (.A(_05070_),
    .B(_05239_),
    .Y(_05243_));
 sky130_fd_sc_hd__o21ai_1 _14282_ (.A1(net115),
    .A2(_05243_),
    .B1(_05242_),
    .Y(_05244_));
 sky130_fd_sc_hd__and2b_1 _14283_ (.A_N(_05244_),
    .B(_05238_),
    .X(_05245_));
 sky130_fd_sc_hd__and2b_1 _14284_ (.A_N(_05238_),
    .B(_05244_),
    .X(_05246_));
 sky130_fd_sc_hd__o31ai_1 _14285_ (.A1(net255),
    .A2(_05245_),
    .A3(_05246_),
    .B1(_05166_),
    .Y(_08663_));
 sky130_fd_sc_hd__mux2_4 _14286_ (.A0(_03352_),
    .A1(_03360_),
    .S(net554),
    .X(_05247_));
 sky130_fd_sc_hd__o21a_1 _14287_ (.A1(_03356_),
    .A2(net204),
    .B1(net205),
    .X(_05248_));
 sky130_fd_sc_hd__a21oi_4 _14288_ (.A1(net539),
    .A2(_05247_),
    .B1(_05248_),
    .Y(_05249_));
 sky130_fd_sc_hd__a22oi_1 _14289_ (.A1(net331),
    .A2(net691),
    .B1(net700),
    .B2(net321),
    .Y(_05250_));
 sky130_fd_sc_hd__and4_1 _14290_ (.A(net321),
    .B(net332),
    .C(net691),
    .D(net700),
    .X(_05252_));
 sky130_fd_sc_hd__or2_1 _14291_ (.A(_05250_),
    .B(_05252_),
    .X(_05253_));
 sky130_fd_sc_hd__nand2_1 _14292_ (.A(net338),
    .B(net682),
    .Y(_05254_));
 sky130_fd_sc_hd__nor2_2 _14293_ (.A(_05253_),
    .B(_05254_),
    .Y(_05255_));
 sky130_fd_sc_hd__and2_1 _14294_ (.A(_05253_),
    .B(_05254_),
    .X(_05256_));
 sky130_fd_sc_hd__nor2_4 _14295_ (.A(_05255_),
    .B(_05256_),
    .Y(_05257_));
 sky130_fd_sc_hd__and2b_1 _14296_ (.A_N(_05172_),
    .B(_05257_),
    .X(_05258_));
 sky130_fd_sc_hd__xor2_4 _14297_ (.A(_05172_),
    .B(_05257_),
    .X(_05259_));
 sky130_fd_sc_hd__o21ba_2 _14298_ (.A1(_05167_),
    .A2(_05170_),
    .B1_N(_05168_),
    .X(_05260_));
 sky130_fd_sc_hd__a22oi_4 _14299_ (.A1(net353),
    .A2(net664),
    .B1(net672),
    .B2(net346),
    .Y(_05261_));
 sky130_fd_sc_hd__nand2_1 _14300_ (.A(net347),
    .B(net664),
    .Y(_05263_));
 sky130_fd_sc_hd__and4_1 _14301_ (.A(net346),
    .B(net353),
    .C(net664),
    .D(net672),
    .X(_05264_));
 sky130_fd_sc_hd__nor2_2 _14302_ (.A(_05261_),
    .B(_05264_),
    .Y(_05265_));
 sky130_fd_sc_hd__nand2_4 _14303_ (.A(net361),
    .B(net656),
    .Y(_05266_));
 sky130_fd_sc_hd__xnor2_4 _14304_ (.A(_05265_),
    .B(_05266_),
    .Y(_05267_));
 sky130_fd_sc_hd__nand2b_2 _14305_ (.A_N(_05260_),
    .B(_05267_),
    .Y(_05268_));
 sky130_fd_sc_hd__xnor2_2 _14306_ (.A(_05260_),
    .B(_05267_),
    .Y(_05269_));
 sky130_fd_sc_hd__o21ba_1 _14307_ (.A1(_05179_),
    .A2(_05182_),
    .B1_N(_05180_),
    .X(_05270_));
 sky130_fd_sc_hd__nand2b_2 _14308_ (.A_N(_05270_),
    .B(_05269_),
    .Y(_05271_));
 sky130_fd_sc_hd__xor2_1 _14309_ (.A(_05269_),
    .B(_05270_),
    .X(_05272_));
 sky130_fd_sc_hd__o21ba_1 _14310_ (.A1(_05185_),
    .A2(_05188_),
    .B1_N(_05184_),
    .X(_05274_));
 sky130_fd_sc_hd__nor2_1 _14311_ (.A(_05272_),
    .B(_05274_),
    .Y(_05275_));
 sky130_fd_sc_hd__and2_1 _14312_ (.A(_05272_),
    .B(_05274_),
    .X(_05276_));
 sky130_fd_sc_hd__or2_1 _14313_ (.A(_05275_),
    .B(_05276_),
    .X(_05277_));
 sky130_fd_sc_hd__or2_2 _14314_ (.A(_05191_),
    .B(_05277_),
    .X(_05278_));
 sky130_fd_sc_hd__nand2_1 _14315_ (.A(_05191_),
    .B(_05277_),
    .Y(_05279_));
 sky130_fd_sc_hd__nand2_1 _14316_ (.A(_05278_),
    .B(_05279_),
    .Y(_05280_));
 sky130_fd_sc_hd__a22oi_1 _14317_ (.A1(net377),
    .A2(net639),
    .B1(net648),
    .B2(net369),
    .Y(_05281_));
 sky130_fd_sc_hd__and4_1 _14318_ (.A(net368),
    .B(net377),
    .C(net639),
    .D(net648),
    .X(_05282_));
 sky130_fd_sc_hd__nor2_1 _14319_ (.A(_05281_),
    .B(_05282_),
    .Y(_05283_));
 sky130_fd_sc_hd__a21oi_1 _14320_ (.A1(net385),
    .A2(net631),
    .B1(_05283_),
    .Y(_05285_));
 sky130_fd_sc_hd__and3_1 _14321_ (.A(net386),
    .B(net630),
    .C(_05283_),
    .X(_05286_));
 sky130_fd_sc_hd__nor2_1 _14322_ (.A(_05285_),
    .B(_05286_),
    .Y(_05287_));
 sky130_fd_sc_hd__o21ba_1 _14323_ (.A1(_05198_),
    .A2(_05201_),
    .B1_N(_05199_),
    .X(_05288_));
 sky130_fd_sc_hd__or3_1 _14324_ (.A(_05285_),
    .B(_05286_),
    .C(_05288_),
    .X(_05289_));
 sky130_fd_sc_hd__xnor2_2 _14325_ (.A(_05287_),
    .B(_05288_),
    .Y(_05290_));
 sky130_fd_sc_hd__nand3_2 _14326_ (.A(net395),
    .B(net622),
    .C(_05290_),
    .Y(_05291_));
 sky130_fd_sc_hd__a21o_1 _14327_ (.A1(net395),
    .A2(net622),
    .B1(_05290_),
    .X(_05292_));
 sky130_fd_sc_hd__nand2_2 _14328_ (.A(_05291_),
    .B(_05292_),
    .Y(_05293_));
 sky130_fd_sc_hd__a21oi_4 _14329_ (.A1(_05204_),
    .A2(_05206_),
    .B1(_05293_),
    .Y(_05294_));
 sky130_fd_sc_hd__and3_1 _14330_ (.A(_05204_),
    .B(_05206_),
    .C(_05293_),
    .X(_05296_));
 sky130_fd_sc_hd__or2_1 _14331_ (.A(_05294_),
    .B(_05296_),
    .X(_05297_));
 sky130_fd_sc_hd__or2_4 _14332_ (.A(_05280_),
    .B(_05297_),
    .X(_05298_));
 sky130_fd_sc_hd__nand2_2 _14333_ (.A(_05280_),
    .B(_05297_),
    .Y(_05299_));
 sky130_fd_sc_hd__o211a_4 _14334_ (.A1(_05194_),
    .A2(_05215_),
    .B1(_05298_),
    .C1(_05299_),
    .X(_05300_));
 sky130_fd_sc_hd__a211oi_4 _14335_ (.A1(_05298_),
    .A2(_05299_),
    .B1(_05194_),
    .C1(_05215_),
    .Y(_05301_));
 sky130_fd_sc_hd__o21a_2 _14336_ (.A1(_05300_),
    .A2(_05301_),
    .B1(_05259_),
    .X(_05302_));
 sky130_fd_sc_hd__nor3_4 _14337_ (.A(_05259_),
    .B(_05300_),
    .C(_05301_),
    .Y(_05303_));
 sky130_fd_sc_hd__a211o_4 _14338_ (.A1(_05176_),
    .A2(_05222_),
    .B1(_05302_),
    .C1(_05303_),
    .X(_05304_));
 sky130_fd_sc_hd__o211ai_4 _14339_ (.A1(_05302_),
    .A2(_05303_),
    .B1(_05176_),
    .C1(_05222_),
    .Y(_05305_));
 sky130_fd_sc_hd__nand3_4 _14340_ (.A(_05218_),
    .B(_05304_),
    .C(_05305_),
    .Y(_05307_));
 sky130_fd_sc_hd__a21o_1 _14341_ (.A1(_05304_),
    .A2(_05305_),
    .B1(_05218_),
    .X(_05308_));
 sky130_fd_sc_hd__and2_1 _14342_ (.A(_05307_),
    .B(_05308_),
    .X(_05309_));
 sky130_fd_sc_hd__o21a_1 _14343_ (.A1(_05225_),
    .A2(_05227_),
    .B1(_05309_),
    .X(_05310_));
 sky130_fd_sc_hd__nor3_1 _14344_ (.A(_05225_),
    .B(_05227_),
    .C(_05309_),
    .Y(_05311_));
 sky130_fd_sc_hd__nor2_1 _14345_ (.A(_05310_),
    .B(_05311_),
    .Y(_05312_));
 sky130_fd_sc_hd__a31oi_4 _14346_ (.A1(net402),
    .A2(net622),
    .A3(_05212_),
    .B1(_05210_),
    .Y(_05313_));
 sky130_fd_sc_hd__and2b_1 _14347_ (.A_N(_05313_),
    .B(_05312_),
    .X(_05314_));
 sky130_fd_sc_hd__xnor2_1 _14348_ (.A(_05312_),
    .B(_05313_),
    .Y(_05315_));
 sky130_fd_sc_hd__o21a_1 _14349_ (.A1(_05229_),
    .A2(_05233_),
    .B1(_05315_),
    .X(_05316_));
 sky130_fd_sc_hd__or3_1 _14350_ (.A(_05229_),
    .B(_05233_),
    .C(_05315_),
    .X(_05318_));
 sky130_fd_sc_hd__and2b_1 _14351_ (.A_N(_05316_),
    .B(_05318_),
    .X(_05319_));
 sky130_fd_sc_hd__or2_1 _14352_ (.A(_05236_),
    .B(_05246_),
    .X(_05320_));
 sky130_fd_sc_hd__nand2_1 _14353_ (.A(_05319_),
    .B(_05320_),
    .Y(_05321_));
 sky130_fd_sc_hd__or2_1 _14354_ (.A(_05319_),
    .B(_05320_),
    .X(_05322_));
 sky130_fd_sc_hd__a31o_1 _14355_ (.A1(net258),
    .A2(_05321_),
    .A3(_05322_),
    .B1(_05249_),
    .X(_08665_));
 sky130_fd_sc_hd__mux2_4 _14356_ (.A0(_03524_),
    .A1(_03527_),
    .S(net554),
    .X(_05323_));
 sky130_fd_sc_hd__o21a_1 _14357_ (.A1(_03521_),
    .A2(net204),
    .B1(net205),
    .X(_05324_));
 sky130_fd_sc_hd__a21oi_4 _14358_ (.A1(net537),
    .A2(_05323_),
    .B1(_05324_),
    .Y(_05325_));
 sky130_fd_sc_hd__a22oi_1 _14359_ (.A1(net332),
    .A2(net681),
    .B1(net691),
    .B2(net321),
    .Y(_05326_));
 sky130_fd_sc_hd__and4_1 _14360_ (.A(net321),
    .B(net332),
    .C(net681),
    .D(net691),
    .X(_05328_));
 sky130_fd_sc_hd__or2_1 _14361_ (.A(_05326_),
    .B(_05328_),
    .X(_05329_));
 sky130_fd_sc_hd__nand2_1 _14362_ (.A(net338),
    .B(net672),
    .Y(_05330_));
 sky130_fd_sc_hd__nor2_1 _14363_ (.A(_05329_),
    .B(_05330_),
    .Y(_05331_));
 sky130_fd_sc_hd__and2_1 _14364_ (.A(_05329_),
    .B(_05330_),
    .X(_05332_));
 sky130_fd_sc_hd__nor2_1 _14365_ (.A(_05331_),
    .B(_05332_),
    .Y(_05333_));
 sky130_fd_sc_hd__nand2_4 _14366_ (.A(net353),
    .B(net657),
    .Y(_05334_));
 sky130_fd_sc_hd__xor2_1 _14367_ (.A(_05263_),
    .B(_05334_),
    .X(_05335_));
 sky130_fd_sc_hd__and3_1 _14368_ (.A(net360),
    .B(net648),
    .C(_05335_),
    .X(_05336_));
 sky130_fd_sc_hd__a21oi_1 _14369_ (.A1(net360),
    .A2(net648),
    .B1(_05335_),
    .Y(_05337_));
 sky130_fd_sc_hd__nor2_1 _14370_ (.A(_05336_),
    .B(_05337_),
    .Y(_05339_));
 sky130_fd_sc_hd__o21ai_2 _14371_ (.A1(_05252_),
    .A2(_05255_),
    .B1(_05339_),
    .Y(_05340_));
 sky130_fd_sc_hd__or3_1 _14372_ (.A(_05252_),
    .B(_05255_),
    .C(_05339_),
    .X(_05341_));
 sky130_fd_sc_hd__and2_2 _14373_ (.A(_05340_),
    .B(_05341_),
    .X(_05342_));
 sky130_fd_sc_hd__o21ba_2 _14374_ (.A1(_05261_),
    .A2(_05266_),
    .B1_N(_05264_),
    .X(_05343_));
 sky130_fd_sc_hd__nand2b_1 _14375_ (.A_N(_05343_),
    .B(_05342_),
    .Y(_05344_));
 sky130_fd_sc_hd__xor2_4 _14376_ (.A(_05342_),
    .B(_05343_),
    .X(_05345_));
 sky130_fd_sc_hd__a21oi_4 _14377_ (.A1(_05268_),
    .A2(_05271_),
    .B1(_05345_),
    .Y(_05346_));
 sky130_fd_sc_hd__and3_1 _14378_ (.A(_05268_),
    .B(_05271_),
    .C(_05345_),
    .X(_05347_));
 sky130_fd_sc_hd__nor2_1 _14379_ (.A(_05346_),
    .B(_05347_),
    .Y(_05348_));
 sky130_fd_sc_hd__and2_2 _14380_ (.A(_05275_),
    .B(_05348_),
    .X(_05350_));
 sky130_fd_sc_hd__nor2_1 _14381_ (.A(_05275_),
    .B(_05348_),
    .Y(_05351_));
 sky130_fd_sc_hd__or2_2 _14382_ (.A(_05350_),
    .B(_05351_),
    .X(_05352_));
 sky130_fd_sc_hd__and2_2 _14383_ (.A(net377),
    .B(net631),
    .X(_05353_));
 sky130_fd_sc_hd__a21oi_2 _14384_ (.A1(net368),
    .A2(net640),
    .B1(_05353_),
    .Y(_05354_));
 sky130_fd_sc_hd__and3_2 _14385_ (.A(net368),
    .B(net640),
    .C(_05353_),
    .X(_05355_));
 sky130_fd_sc_hd__nor2_4 _14386_ (.A(_05354_),
    .B(_05355_),
    .Y(_05356_));
 sky130_fd_sc_hd__nand2_2 _14387_ (.A(net386),
    .B(net622),
    .Y(_05357_));
 sky130_fd_sc_hd__xnor2_4 _14388_ (.A(_05356_),
    .B(_05357_),
    .Y(_05358_));
 sky130_fd_sc_hd__or2_4 _14389_ (.A(_05282_),
    .B(_05286_),
    .X(_05359_));
 sky130_fd_sc_hd__xnor2_2 _14390_ (.A(_05358_),
    .B(_05359_),
    .Y(_05361_));
 sky130_fd_sc_hd__a21oi_2 _14391_ (.A1(_05289_),
    .A2(_05291_),
    .B1(_05361_),
    .Y(_05362_));
 sky130_fd_sc_hd__inv_2 _14392_ (.A(_05362_),
    .Y(_05363_));
 sky130_fd_sc_hd__and3_1 _14393_ (.A(_05289_),
    .B(_05291_),
    .C(_05361_),
    .X(_05364_));
 sky130_fd_sc_hd__or2_2 _14394_ (.A(_05362_),
    .B(_05364_),
    .X(_05365_));
 sky130_fd_sc_hd__nor2_4 _14395_ (.A(_05352_),
    .B(_05365_),
    .Y(_05366_));
 sky130_fd_sc_hd__and2_1 _14396_ (.A(_05352_),
    .B(_05365_),
    .X(_05367_));
 sky130_fd_sc_hd__a211o_1 _14397_ (.A1(_05278_),
    .A2(_05298_),
    .B1(_05366_),
    .C1(_05367_),
    .X(_05368_));
 sky130_fd_sc_hd__o211ai_2 _14398_ (.A1(_05366_),
    .A2(_05367_),
    .B1(_05278_),
    .C1(_05298_),
    .Y(_05369_));
 sky130_fd_sc_hd__a21o_1 _14399_ (.A1(_05368_),
    .A2(_05369_),
    .B1(_05333_),
    .X(_05370_));
 sky130_fd_sc_hd__and3_1 _14400_ (.A(_05333_),
    .B(_05368_),
    .C(_05369_),
    .X(_05372_));
 sky130_fd_sc_hd__inv_2 _14401_ (.A(_05372_),
    .Y(_05373_));
 sky130_fd_sc_hd__o211a_1 _14402_ (.A1(_05258_),
    .A2(_05303_),
    .B1(_05370_),
    .C1(_05373_),
    .X(_05374_));
 sky130_fd_sc_hd__inv_2 _14403_ (.A(_05374_),
    .Y(_05375_));
 sky130_fd_sc_hd__a211o_2 _14404_ (.A1(_05370_),
    .A2(_05373_),
    .B1(_05258_),
    .C1(_05303_),
    .X(_05376_));
 sky130_fd_sc_hd__and3_4 _14405_ (.A(_05300_),
    .B(_05375_),
    .C(_05376_),
    .X(_05377_));
 sky130_fd_sc_hd__a21oi_4 _14406_ (.A1(_05375_),
    .A2(_05376_),
    .B1(_05300_),
    .Y(_05378_));
 sky130_fd_sc_hd__a211o_4 _14407_ (.A1(_05304_),
    .A2(_05307_),
    .B1(_05377_),
    .C1(_05378_),
    .X(_05379_));
 sky130_fd_sc_hd__o211ai_4 _14408_ (.A1(_05377_),
    .A2(_05378_),
    .B1(_05304_),
    .C1(_05307_),
    .Y(_05380_));
 sky130_fd_sc_hd__nand3_4 _14409_ (.A(_05294_),
    .B(_05379_),
    .C(_05380_),
    .Y(_05381_));
 sky130_fd_sc_hd__a21o_1 _14410_ (.A1(_05379_),
    .A2(_05380_),
    .B1(_05294_),
    .X(_05383_));
 sky130_fd_sc_hd__and2_1 _14411_ (.A(_05381_),
    .B(_05383_),
    .X(_05384_));
 sky130_fd_sc_hd__o21a_2 _14412_ (.A1(_05310_),
    .A2(_05314_),
    .B1(_05384_),
    .X(_05385_));
 sky130_fd_sc_hd__nor3_1 _14413_ (.A(_05310_),
    .B(_05314_),
    .C(_05384_),
    .Y(_05386_));
 sky130_fd_sc_hd__nor2_1 _14414_ (.A(_05385_),
    .B(_05386_),
    .Y(_05387_));
 sky130_fd_sc_hd__o21a_1 _14415_ (.A1(_05236_),
    .A2(_05316_),
    .B1(_05318_),
    .X(_05388_));
 sky130_fd_sc_hd__and2b_1 _14416_ (.A_N(_05238_),
    .B(_05319_),
    .X(_05389_));
 sky130_fd_sc_hd__a21o_1 _14417_ (.A1(_05244_),
    .A2(_05389_),
    .B1(_05388_),
    .X(_05390_));
 sky130_fd_sc_hd__or2_1 _14418_ (.A(_05387_),
    .B(_05390_),
    .X(_05391_));
 sky130_fd_sc_hd__nand2_1 _14419_ (.A(_05387_),
    .B(_05390_),
    .Y(_05392_));
 sky130_fd_sc_hd__a31o_1 _14420_ (.A1(net258),
    .A2(_05391_),
    .A3(_05392_),
    .B1(_05325_),
    .X(_08666_));
 sky130_fd_sc_hd__mux2_4 _14421_ (.A0(_03677_),
    .A1(_03684_),
    .S(net553),
    .X(_05394_));
 sky130_fd_sc_hd__o21a_1 _14422_ (.A1(_03680_),
    .A2(net204),
    .B1(net205),
    .X(_05395_));
 sky130_fd_sc_hd__a21oi_4 _14423_ (.A1(net537),
    .A2(_05394_),
    .B1(_05395_),
    .Y(_05396_));
 sky130_fd_sc_hd__nor2_2 _14424_ (.A(_05374_),
    .B(_05377_),
    .Y(_05397_));
 sky130_fd_sc_hd__a22oi_1 _14425_ (.A1(net332),
    .A2(net672),
    .B1(net681),
    .B2(net321),
    .Y(_05398_));
 sky130_fd_sc_hd__and4_1 _14426_ (.A(net321),
    .B(net332),
    .C(net672),
    .D(net681),
    .X(_05399_));
 sky130_fd_sc_hd__or2_1 _14427_ (.A(_05398_),
    .B(_05399_),
    .X(_05400_));
 sky130_fd_sc_hd__nand2_1 _14428_ (.A(net339),
    .B(net665),
    .Y(_05401_));
 sky130_fd_sc_hd__nor2_1 _14429_ (.A(_05400_),
    .B(_05401_),
    .Y(_05402_));
 sky130_fd_sc_hd__and2_1 _14430_ (.A(_05400_),
    .B(_05401_),
    .X(_05404_));
 sky130_fd_sc_hd__nor2_1 _14431_ (.A(_05402_),
    .B(_05404_),
    .Y(_05405_));
 sky130_fd_sc_hd__a22o_1 _14432_ (.A1(net353),
    .A2(net649),
    .B1(net656),
    .B2(net347),
    .X(_05406_));
 sky130_fd_sc_hd__nand2_8 _14433_ (.A(net343),
    .B(net649),
    .Y(_05407_));
 sky130_fd_sc_hd__inv_2 _14434_ (.A(_05407_),
    .Y(_05408_));
 sky130_fd_sc_hd__o21a_1 _14435_ (.A1(_05334_),
    .A2(_05407_),
    .B1(_05406_),
    .X(_05409_));
 sky130_fd_sc_hd__a21oi_1 _14436_ (.A1(net360),
    .A2(net639),
    .B1(_05409_),
    .Y(_05410_));
 sky130_fd_sc_hd__and3_1 _14437_ (.A(net360),
    .B(net639),
    .C(_05409_),
    .X(_05411_));
 sky130_fd_sc_hd__nor2_1 _14438_ (.A(_05410_),
    .B(_05411_),
    .Y(_05412_));
 sky130_fd_sc_hd__o21a_1 _14439_ (.A1(_05328_),
    .A2(_05331_),
    .B1(_05412_),
    .X(_05413_));
 sky130_fd_sc_hd__nor3_1 _14440_ (.A(_05328_),
    .B(_05331_),
    .C(_05412_),
    .Y(_05415_));
 sky130_fd_sc_hd__nor2_1 _14441_ (.A(_05413_),
    .B(_05415_),
    .Y(_05416_));
 sky130_fd_sc_hd__o21ba_2 _14442_ (.A1(_05263_),
    .A2(_05334_),
    .B1_N(_05336_),
    .X(_05417_));
 sky130_fd_sc_hd__xor2_2 _14443_ (.A(_05416_),
    .B(_05417_),
    .X(_05418_));
 sky130_fd_sc_hd__a21o_2 _14444_ (.A1(_05340_),
    .A2(_05344_),
    .B1(_05418_),
    .X(_05419_));
 sky130_fd_sc_hd__nand3_2 _14445_ (.A(_05340_),
    .B(_05344_),
    .C(_05418_),
    .Y(_05420_));
 sky130_fd_sc_hd__nand3_4 _14446_ (.A(_05346_),
    .B(_05419_),
    .C(_05420_),
    .Y(_05421_));
 sky130_fd_sc_hd__a21o_1 _14447_ (.A1(_05419_),
    .A2(_05420_),
    .B1(_05346_),
    .X(_05422_));
 sky130_fd_sc_hd__a22oi_1 _14448_ (.A1(net378),
    .A2(net622),
    .B1(net631),
    .B2(net368),
    .Y(_05423_));
 sky130_fd_sc_hd__nand2_1 _14449_ (.A(net368),
    .B(net622),
    .Y(_05424_));
 sky130_fd_sc_hd__and3_2 _14450_ (.A(net368),
    .B(net622),
    .C(_05353_),
    .X(_05426_));
 sky130_fd_sc_hd__nor2_1 _14451_ (.A(_05423_),
    .B(_05426_),
    .Y(_05427_));
 sky130_fd_sc_hd__a31o_1 _14452_ (.A1(net385),
    .A2(net622),
    .A3(_05356_),
    .B1(_05355_),
    .X(_05428_));
 sky130_fd_sc_hd__nand2_1 _14453_ (.A(_05427_),
    .B(_05428_),
    .Y(_05429_));
 sky130_fd_sc_hd__or2_1 _14454_ (.A(_05427_),
    .B(_05428_),
    .X(_05430_));
 sky130_fd_sc_hd__and2_1 _14455_ (.A(_05429_),
    .B(_05430_),
    .X(_05431_));
 sky130_fd_sc_hd__nand3_2 _14456_ (.A(_05358_),
    .B(_05359_),
    .C(_05431_),
    .Y(_05432_));
 sky130_fd_sc_hd__a21o_1 _14457_ (.A1(_05358_),
    .A2(_05359_),
    .B1(_05431_),
    .X(_05433_));
 sky130_fd_sc_hd__and2_2 _14458_ (.A(_05432_),
    .B(_05433_),
    .X(_05434_));
 sky130_fd_sc_hd__nand3_4 _14459_ (.A(_05421_),
    .B(_05422_),
    .C(_05434_),
    .Y(_05435_));
 sky130_fd_sc_hd__a21o_1 _14460_ (.A1(_05421_),
    .A2(_05422_),
    .B1(_05434_),
    .X(_05437_));
 sky130_fd_sc_hd__o211ai_4 _14461_ (.A1(_05350_),
    .A2(_05366_),
    .B1(_05435_),
    .C1(_05437_),
    .Y(_05438_));
 sky130_fd_sc_hd__a211o_1 _14462_ (.A1(_05435_),
    .A2(_05437_),
    .B1(_05350_),
    .C1(_05366_),
    .X(_05439_));
 sky130_fd_sc_hd__nand3_2 _14463_ (.A(_05405_),
    .B(_05438_),
    .C(_05439_),
    .Y(_05440_));
 sky130_fd_sc_hd__a21o_1 _14464_ (.A1(_05438_),
    .A2(_05439_),
    .B1(_05405_),
    .X(_05441_));
 sky130_fd_sc_hd__nand2_2 _14465_ (.A(_05440_),
    .B(_05441_),
    .Y(_05442_));
 sky130_fd_sc_hd__and2_2 _14466_ (.A(_05368_),
    .B(_05373_),
    .X(_05443_));
 sky130_fd_sc_hd__xnor2_2 _14467_ (.A(_05442_),
    .B(_05443_),
    .Y(_05444_));
 sky130_fd_sc_hd__nor2_1 _14468_ (.A(_05397_),
    .B(_05444_),
    .Y(_05445_));
 sky130_fd_sc_hd__xnor2_1 _14469_ (.A(_05397_),
    .B(_05444_),
    .Y(_05446_));
 sky130_fd_sc_hd__nor2_1 _14470_ (.A(_05363_),
    .B(_05446_),
    .Y(_05448_));
 sky130_fd_sc_hd__and2_1 _14471_ (.A(_05363_),
    .B(_05446_),
    .X(_05449_));
 sky130_fd_sc_hd__or2_2 _14472_ (.A(_05448_),
    .B(_05449_),
    .X(_05450_));
 sky130_fd_sc_hd__nand3_2 _14473_ (.A(_05379_),
    .B(_05381_),
    .C(_05450_),
    .Y(_05451_));
 sky130_fd_sc_hd__a21oi_2 _14474_ (.A1(_05379_),
    .A2(_05381_),
    .B1(_05450_),
    .Y(_05452_));
 sky130_fd_sc_hd__inv_2 _14475_ (.A(_05452_),
    .Y(_05453_));
 sky130_fd_sc_hd__nand2_1 _14476_ (.A(_05451_),
    .B(_05453_),
    .Y(_05454_));
 sky130_fd_sc_hd__a21oi_1 _14477_ (.A1(_05387_),
    .A2(_05390_),
    .B1(_05385_),
    .Y(_05455_));
 sky130_fd_sc_hd__or2_1 _14478_ (.A(_05454_),
    .B(_05455_),
    .X(_05456_));
 sky130_fd_sc_hd__nand2_1 _14479_ (.A(_05454_),
    .B(_05455_),
    .Y(_05457_));
 sky130_fd_sc_hd__a31o_1 _14480_ (.A1(net261),
    .A2(_05456_),
    .A3(_05457_),
    .B1(_05396_),
    .X(_08667_));
 sky130_fd_sc_hd__mux2_4 _14481_ (.A0(_03690_),
    .A1(_03695_),
    .S(net308),
    .X(_05459_));
 sky130_fd_sc_hd__o31a_1 _14482_ (.A1(net300),
    .A2(_03697_),
    .A3(net204),
    .B1(net205),
    .X(_05460_));
 sky130_fd_sc_hd__a21oi_4 _14483_ (.A1(net537),
    .A2(_05459_),
    .B1(_05460_),
    .Y(_05461_));
 sky130_fd_sc_hd__a22oi_1 _14484_ (.A1(net330),
    .A2(net664),
    .B1(net672),
    .B2(net320),
    .Y(_05462_));
 sky130_fd_sc_hd__and4_1 _14485_ (.A(net320),
    .B(net329),
    .C(net665),
    .D(net672),
    .X(_05463_));
 sky130_fd_sc_hd__or2_1 _14486_ (.A(_05462_),
    .B(_05463_),
    .X(_05464_));
 sky130_fd_sc_hd__nand2_1 _14487_ (.A(net337),
    .B(net657),
    .Y(_05465_));
 sky130_fd_sc_hd__nor2_1 _14488_ (.A(_05464_),
    .B(_05465_),
    .Y(_05466_));
 sky130_fd_sc_hd__and2_1 _14489_ (.A(_05464_),
    .B(_05465_),
    .X(_05467_));
 sky130_fd_sc_hd__nor2_1 _14490_ (.A(_05466_),
    .B(_05467_),
    .Y(_05469_));
 sky130_fd_sc_hd__nand2_1 _14491_ (.A(net353),
    .B(net638),
    .Y(_05470_));
 sky130_fd_sc_hd__xor2_1 _14492_ (.A(_05407_),
    .B(_05470_),
    .X(_05471_));
 sky130_fd_sc_hd__and3_1 _14493_ (.A(net360),
    .B(net629),
    .C(_05471_),
    .X(_05472_));
 sky130_fd_sc_hd__a21oi_1 _14494_ (.A1(net360),
    .A2(net629),
    .B1(_05471_),
    .Y(_05473_));
 sky130_fd_sc_hd__nor2_1 _14495_ (.A(_05472_),
    .B(_05473_),
    .Y(_05474_));
 sky130_fd_sc_hd__o21ai_2 _14496_ (.A1(_05399_),
    .A2(_05402_),
    .B1(_05474_),
    .Y(_05475_));
 sky130_fd_sc_hd__or3_1 _14497_ (.A(_05399_),
    .B(_05402_),
    .C(_05474_),
    .X(_05476_));
 sky130_fd_sc_hd__and2_1 _14498_ (.A(_05475_),
    .B(_05476_),
    .X(_05477_));
 sky130_fd_sc_hd__o21ba_1 _14499_ (.A1(_05334_),
    .A2(_05407_),
    .B1_N(_05411_),
    .X(_05478_));
 sky130_fd_sc_hd__nand2b_1 _14500_ (.A_N(_05477_),
    .B(_05478_),
    .Y(_05480_));
 sky130_fd_sc_hd__nand2b_1 _14501_ (.A_N(_05478_),
    .B(_05477_),
    .Y(_05481_));
 sky130_fd_sc_hd__nand2_1 _14502_ (.A(_05480_),
    .B(_05481_),
    .Y(_05482_));
 sky130_fd_sc_hd__o21ba_1 _14503_ (.A1(_05415_),
    .A2(_05417_),
    .B1_N(_05413_),
    .X(_05483_));
 sky130_fd_sc_hd__nor2_1 _14504_ (.A(_05482_),
    .B(_05483_),
    .Y(_05484_));
 sky130_fd_sc_hd__and2_1 _14505_ (.A(_05482_),
    .B(_05483_),
    .X(_05485_));
 sky130_fd_sc_hd__nor2_1 _14506_ (.A(_05484_),
    .B(_05485_),
    .Y(_05486_));
 sky130_fd_sc_hd__nand2b_1 _14507_ (.A_N(_05419_),
    .B(_05486_),
    .Y(_05487_));
 sky130_fd_sc_hd__xnor2_1 _14508_ (.A(_05419_),
    .B(_05486_),
    .Y(_05488_));
 sky130_fd_sc_hd__nor3_2 _14509_ (.A(_05353_),
    .B(_05424_),
    .C(_05429_),
    .Y(_05489_));
 sky130_fd_sc_hd__inv_2 _14510_ (.A(_05489_),
    .Y(_05491_));
 sky130_fd_sc_hd__o21a_1 _14511_ (.A1(_05353_),
    .A2(_05424_),
    .B1(_05429_),
    .X(_05492_));
 sky130_fd_sc_hd__nor2_1 _14512_ (.A(_05489_),
    .B(_05492_),
    .Y(_05493_));
 sky130_fd_sc_hd__nand2_1 _14513_ (.A(_05488_),
    .B(_05493_),
    .Y(_05494_));
 sky130_fd_sc_hd__or2_1 _14514_ (.A(_05488_),
    .B(_05493_),
    .X(_05495_));
 sky130_fd_sc_hd__nand2_1 _14515_ (.A(_05494_),
    .B(_05495_),
    .Y(_05496_));
 sky130_fd_sc_hd__a21o_1 _14516_ (.A1(_05421_),
    .A2(_05435_),
    .B1(_05496_),
    .X(_05497_));
 sky130_fd_sc_hd__clkinv_2 _14517_ (.A(_05497_),
    .Y(_05498_));
 sky130_fd_sc_hd__nand3_1 _14518_ (.A(_05421_),
    .B(_05435_),
    .C(_05496_),
    .Y(_05499_));
 sky130_fd_sc_hd__and3_4 _14519_ (.A(_05469_),
    .B(_05497_),
    .C(_05499_),
    .X(_05500_));
 sky130_fd_sc_hd__a21oi_1 _14520_ (.A1(_05497_),
    .A2(_05499_),
    .B1(_05469_),
    .Y(_05502_));
 sky130_fd_sc_hd__a211o_2 _14521_ (.A1(_05438_),
    .A2(_05440_),
    .B1(_05500_),
    .C1(_05502_),
    .X(_05503_));
 sky130_fd_sc_hd__o211ai_1 _14522_ (.A1(_05500_),
    .A2(_05502_),
    .B1(_05438_),
    .C1(_05440_),
    .Y(_05504_));
 sky130_fd_sc_hd__nand2_1 _14523_ (.A(_05503_),
    .B(_05504_),
    .Y(_05505_));
 sky130_fd_sc_hd__or3_2 _14524_ (.A(_05442_),
    .B(_05443_),
    .C(_05505_),
    .X(_05506_));
 sky130_fd_sc_hd__o21ai_1 _14525_ (.A1(_05442_),
    .A2(_05443_),
    .B1(_05505_),
    .Y(_05507_));
 sky130_fd_sc_hd__nand2_1 _14526_ (.A(_05506_),
    .B(_05507_),
    .Y(_05508_));
 sky130_fd_sc_hd__or2_1 _14527_ (.A(_05432_),
    .B(_05508_),
    .X(_05509_));
 sky130_fd_sc_hd__nand2_1 _14528_ (.A(_05432_),
    .B(_05508_),
    .Y(_05510_));
 sky130_fd_sc_hd__and2_1 _14529_ (.A(_05509_),
    .B(_05510_),
    .X(_05511_));
 sky130_fd_sc_hd__o21ai_2 _14530_ (.A1(_05445_),
    .A2(_05448_),
    .B1(_05511_),
    .Y(_05513_));
 sky130_fd_sc_hd__or3_1 _14531_ (.A(_05445_),
    .B(_05448_),
    .C(_05511_),
    .X(_05514_));
 sky130_fd_sc_hd__and2_1 _14532_ (.A(_05513_),
    .B(_05514_),
    .X(_05515_));
 sky130_fd_sc_hd__and3_1 _14533_ (.A(_05387_),
    .B(_05451_),
    .C(_05453_),
    .X(_05516_));
 sky130_fd_sc_hd__nand2_2 _14534_ (.A(_05389_),
    .B(_05516_),
    .Y(_05517_));
 sky130_fd_sc_hd__o21ai_2 _14535_ (.A1(_05385_),
    .A2(_05452_),
    .B1(_05451_),
    .Y(_05518_));
 sky130_fd_sc_hd__o2bb2a_1 _14536_ (.A1_N(_05388_),
    .A2_N(_05516_),
    .B1(_05517_),
    .B2(_05242_),
    .X(_05519_));
 sky130_fd_sc_hd__o311ai_4 _14537_ (.A1(net115),
    .A2(_05243_),
    .A3(_05517_),
    .B1(_05518_),
    .C1(_05519_),
    .Y(_05520_));
 sky130_fd_sc_hd__or2_1 _14538_ (.A(_05515_),
    .B(_05520_),
    .X(_05521_));
 sky130_fd_sc_hd__nand2_1 _14539_ (.A(_05515_),
    .B(_05520_),
    .Y(_05522_));
 sky130_fd_sc_hd__a31o_1 _14540_ (.A1(net258),
    .A2(_05521_),
    .A3(_05522_),
    .B1(_05461_),
    .X(_08668_));
 sky130_fd_sc_hd__a31o_2 _14541_ (.A1(net554),
    .A2(net570),
    .A3(_02614_),
    .B1(net537),
    .X(_05524_));
 sky130_fd_sc_hd__o22a_2 _14542_ (.A1(net206),
    .A2(_03860_),
    .B1(net204),
    .B2(_03858_),
    .X(_05525_));
 sky130_fd_sc_hd__nand2_2 _14543_ (.A(net208),
    .B(_05525_),
    .Y(_05526_));
 sky130_fd_sc_hd__a22oi_4 _14544_ (.A1(net329),
    .A2(net658),
    .B1(net666),
    .B2(net319),
    .Y(_05527_));
 sky130_fd_sc_hd__and4_2 _14545_ (.A(net319),
    .B(net329),
    .C(net658),
    .D(net666),
    .X(_05528_));
 sky130_fd_sc_hd__nand2_1 _14546_ (.A(net336),
    .B(net647),
    .Y(_05529_));
 sky130_fd_sc_hd__o21a_1 _14547_ (.A1(_05527_),
    .A2(_05528_),
    .B1(_05529_),
    .X(_05530_));
 sky130_fd_sc_hd__nor3_2 _14548_ (.A(_05527_),
    .B(_05528_),
    .C(_05529_),
    .Y(_05531_));
 sky130_fd_sc_hd__nor2_2 _14549_ (.A(_05530_),
    .B(_05531_),
    .Y(_05532_));
 sky130_fd_sc_hd__nand2_1 _14550_ (.A(net354),
    .B(net629),
    .Y(_05534_));
 sky130_fd_sc_hd__a21boi_1 _14551_ (.A1(net343),
    .A2(net637),
    .B1_N(_05534_),
    .Y(_05535_));
 sky130_fd_sc_hd__and4_1 _14552_ (.A(net343),
    .B(net354),
    .C(net629),
    .D(net637),
    .X(_05536_));
 sky130_fd_sc_hd__nor2_1 _14553_ (.A(_05535_),
    .B(_05536_),
    .Y(_05537_));
 sky130_fd_sc_hd__nand2_1 _14554_ (.A(net361),
    .B(net620),
    .Y(_05538_));
 sky130_fd_sc_hd__xnor2_1 _14555_ (.A(_05537_),
    .B(_05538_),
    .Y(_05539_));
 sky130_fd_sc_hd__o21a_1 _14556_ (.A1(_05463_),
    .A2(_05466_),
    .B1(_05539_),
    .X(_05540_));
 sky130_fd_sc_hd__nor3_1 _14557_ (.A(_05463_),
    .B(_05466_),
    .C(_05539_),
    .Y(_05541_));
 sky130_fd_sc_hd__nor2_1 _14558_ (.A(_05540_),
    .B(_05541_),
    .Y(_05542_));
 sky130_fd_sc_hd__o21ba_2 _14559_ (.A1(_05407_),
    .A2(_05470_),
    .B1_N(_05472_),
    .X(_05543_));
 sky130_fd_sc_hd__xor2_2 _14560_ (.A(_05542_),
    .B(_05543_),
    .X(_05545_));
 sky130_fd_sc_hd__a21o_2 _14561_ (.A1(_05475_),
    .A2(_05481_),
    .B1(_05545_),
    .X(_05546_));
 sky130_fd_sc_hd__nand3_1 _14562_ (.A(_05475_),
    .B(_05481_),
    .C(_05545_),
    .Y(_05547_));
 sky130_fd_sc_hd__and2_1 _14563_ (.A(_05546_),
    .B(_05547_),
    .X(_05548_));
 sky130_fd_sc_hd__and3_1 _14564_ (.A(_05484_),
    .B(_05546_),
    .C(_05547_),
    .X(_05549_));
 sky130_fd_sc_hd__nor2_1 _14565_ (.A(_05484_),
    .B(_05548_),
    .Y(_05550_));
 sky130_fd_sc_hd__nor2_2 _14566_ (.A(_05549_),
    .B(_05550_),
    .Y(_05551_));
 sky130_fd_sc_hd__xnor2_2 _14567_ (.A(_05426_),
    .B(_05551_),
    .Y(_05552_));
 sky130_fd_sc_hd__a21o_2 _14568_ (.A1(_05487_),
    .A2(_05494_),
    .B1(_05552_),
    .X(_05553_));
 sky130_fd_sc_hd__nand3_2 _14569_ (.A(_05487_),
    .B(_05494_),
    .C(_05552_),
    .Y(_05554_));
 sky130_fd_sc_hd__nand3_4 _14570_ (.A(_05532_),
    .B(_05553_),
    .C(_05554_),
    .Y(_05556_));
 sky130_fd_sc_hd__a21o_2 _14571_ (.A1(_05553_),
    .A2(_05554_),
    .B1(_05532_),
    .X(_05557_));
 sky130_fd_sc_hd__o211ai_4 _14572_ (.A1(_05498_),
    .A2(_05500_),
    .B1(_05556_),
    .C1(_05557_),
    .Y(_05558_));
 sky130_fd_sc_hd__a211oi_2 _14573_ (.A1(_05556_),
    .A2(_05557_),
    .B1(_05498_),
    .C1(_05500_),
    .Y(_05559_));
 sky130_fd_sc_hd__inv_2 _14574_ (.A(_05559_),
    .Y(_05560_));
 sky130_fd_sc_hd__nand2_1 _14575_ (.A(_05558_),
    .B(_05560_),
    .Y(_05561_));
 sky130_fd_sc_hd__nor2_1 _14576_ (.A(_05503_),
    .B(_05561_),
    .Y(_05562_));
 sky130_fd_sc_hd__xnor2_1 _14577_ (.A(_05503_),
    .B(_05561_),
    .Y(_05563_));
 sky130_fd_sc_hd__nor2_1 _14578_ (.A(_05491_),
    .B(_05563_),
    .Y(_05564_));
 sky130_fd_sc_hd__and2_1 _14579_ (.A(_05491_),
    .B(_05563_),
    .X(_05565_));
 sky130_fd_sc_hd__or2_1 _14580_ (.A(_05564_),
    .B(_05565_),
    .X(_05567_));
 sky130_fd_sc_hd__a21o_1 _14581_ (.A1(_05506_),
    .A2(_05509_),
    .B1(_05567_),
    .X(_05568_));
 sky130_fd_sc_hd__inv_2 _14582_ (.A(_05568_),
    .Y(_05569_));
 sky130_fd_sc_hd__and3_1 _14583_ (.A(_05506_),
    .B(_05509_),
    .C(_05567_),
    .X(_05570_));
 sky130_fd_sc_hd__nor2_1 _14584_ (.A(_05569_),
    .B(_05570_),
    .Y(_05571_));
 sky130_fd_sc_hd__nand2_1 _14585_ (.A(_05513_),
    .B(_05522_),
    .Y(_05572_));
 sky130_fd_sc_hd__or2_1 _14586_ (.A(_05571_),
    .B(_05572_),
    .X(_05573_));
 sky130_fd_sc_hd__nand2_1 _14587_ (.A(_05571_),
    .B(_05572_),
    .Y(_05574_));
 sky130_fd_sc_hd__a32o_1 _14588_ (.A1(net258),
    .A2(_05573_),
    .A3(_05574_),
    .B1(_05524_),
    .B2(_05526_),
    .X(_08669_));
 sky130_fd_sc_hd__mux2_2 _14589_ (.A0(_04000_),
    .A1(_04002_),
    .S(net309),
    .X(_05575_));
 sky130_fd_sc_hd__nand2_1 _14590_ (.A(net538),
    .B(_05575_),
    .Y(_05577_));
 sky130_fd_sc_hd__a31o_1 _14591_ (.A1(net568),
    .A2(_02830_),
    .A3(_04527_),
    .B1(_03685_),
    .X(_05578_));
 sky130_fd_sc_hd__a22oi_4 _14592_ (.A1(net329),
    .A2(net646),
    .B1(net658),
    .B2(net319),
    .Y(_05579_));
 sky130_fd_sc_hd__and4_1 _14593_ (.A(net319),
    .B(net329),
    .C(net646),
    .D(net658),
    .X(_05580_));
 sky130_fd_sc_hd__or2_2 _14594_ (.A(_05579_),
    .B(_05580_),
    .X(_05581_));
 sky130_fd_sc_hd__and2_4 _14595_ (.A(net336),
    .B(net637),
    .X(_05582_));
 sky130_fd_sc_hd__nand2_2 _14596_ (.A(net336),
    .B(net637),
    .Y(_05583_));
 sky130_fd_sc_hd__xnor2_2 _14597_ (.A(_05581_),
    .B(_05582_),
    .Y(_05584_));
 sky130_fd_sc_hd__a22oi_1 _14598_ (.A1(net354),
    .A2(net621),
    .B1(net629),
    .B2(net343),
    .Y(_05585_));
 sky130_fd_sc_hd__and4_1 _14599_ (.A(net343),
    .B(net354),
    .C(net621),
    .D(net629),
    .X(_05586_));
 sky130_fd_sc_hd__nor2_1 _14600_ (.A(_05585_),
    .B(_05586_),
    .Y(_05588_));
 sky130_fd_sc_hd__or3_1 _14601_ (.A(_05528_),
    .B(_05531_),
    .C(_05588_),
    .X(_05589_));
 sky130_fd_sc_hd__o21ai_2 _14602_ (.A1(_05528_),
    .A2(_05531_),
    .B1(_05588_),
    .Y(_05590_));
 sky130_fd_sc_hd__and2_1 _14603_ (.A(_05589_),
    .B(_05590_),
    .X(_05591_));
 sky130_fd_sc_hd__o21ba_1 _14604_ (.A1(_05535_),
    .A2(_05538_),
    .B1_N(_05536_),
    .X(_05592_));
 sky130_fd_sc_hd__nand2b_1 _14605_ (.A_N(_05592_),
    .B(_05591_),
    .Y(_05593_));
 sky130_fd_sc_hd__xor2_1 _14606_ (.A(_05591_),
    .B(_05592_),
    .X(_05594_));
 sky130_fd_sc_hd__o21ba_1 _14607_ (.A1(_05541_),
    .A2(_05543_),
    .B1_N(_05540_),
    .X(_05595_));
 sky130_fd_sc_hd__nor2_1 _14608_ (.A(_05594_),
    .B(_05595_),
    .Y(_05596_));
 sky130_fd_sc_hd__and2_1 _14609_ (.A(_05594_),
    .B(_05595_),
    .X(_05597_));
 sky130_fd_sc_hd__nor2_1 _14610_ (.A(_05596_),
    .B(_05597_),
    .Y(_05599_));
 sky130_fd_sc_hd__and2b_1 _14611_ (.A_N(_05546_),
    .B(_05599_),
    .X(_05600_));
 sky130_fd_sc_hd__xnor2_1 _14612_ (.A(_05546_),
    .B(_05599_),
    .Y(_05601_));
 sky130_fd_sc_hd__a21oi_1 _14613_ (.A1(_05426_),
    .A2(_05551_),
    .B1(_05549_),
    .Y(_05602_));
 sky130_fd_sc_hd__and2b_1 _14614_ (.A_N(_05602_),
    .B(_05601_),
    .X(_05603_));
 sky130_fd_sc_hd__and2b_1 _14615_ (.A_N(_05601_),
    .B(_05602_),
    .X(_05604_));
 sky130_fd_sc_hd__nor2_1 _14616_ (.A(_05603_),
    .B(_05604_),
    .Y(_05605_));
 sky130_fd_sc_hd__and2_1 _14617_ (.A(_05584_),
    .B(_05605_),
    .X(_05606_));
 sky130_fd_sc_hd__nor2_1 _14618_ (.A(_05584_),
    .B(_05605_),
    .Y(_05607_));
 sky130_fd_sc_hd__or2_1 _14619_ (.A(_05606_),
    .B(_05607_),
    .X(_05608_));
 sky130_fd_sc_hd__a21oi_2 _14620_ (.A1(_05553_),
    .A2(_05556_),
    .B1(_05608_),
    .Y(_05610_));
 sky130_fd_sc_hd__and3_1 _14621_ (.A(_05553_),
    .B(_05556_),
    .C(_05608_),
    .X(_05611_));
 sky130_fd_sc_hd__or2_1 _14622_ (.A(_05610_),
    .B(_05611_),
    .X(_05612_));
 sky130_fd_sc_hd__nor2_2 _14623_ (.A(_05558_),
    .B(_05612_),
    .Y(_05613_));
 sky130_fd_sc_hd__and2_1 _14624_ (.A(_05558_),
    .B(_05612_),
    .X(_05614_));
 sky130_fd_sc_hd__nor2_1 _14625_ (.A(_05613_),
    .B(_05614_),
    .Y(_05615_));
 sky130_fd_sc_hd__o21ai_2 _14626_ (.A1(_05562_),
    .A2(_05564_),
    .B1(_05615_),
    .Y(_05616_));
 sky130_fd_sc_hd__or3_1 _14627_ (.A(_05562_),
    .B(_05564_),
    .C(_05615_),
    .X(_05617_));
 sky130_fd_sc_hd__and2_2 _14628_ (.A(_05616_),
    .B(_05617_),
    .X(_05618_));
 sky130_fd_sc_hd__and3_2 _14629_ (.A(_05515_),
    .B(_05520_),
    .C(_05571_),
    .X(_05619_));
 sky130_fd_sc_hd__a21oi_1 _14630_ (.A1(_05513_),
    .A2(_05568_),
    .B1(_05570_),
    .Y(_05621_));
 sky130_fd_sc_hd__or2_1 _14631_ (.A(_05619_),
    .B(_05621_),
    .X(_05622_));
 sky130_fd_sc_hd__or2_1 _14632_ (.A(_05618_),
    .B(_05622_),
    .X(_05623_));
 sky130_fd_sc_hd__nand2_1 _14633_ (.A(_05618_),
    .B(_05622_),
    .Y(_05624_));
 sky130_fd_sc_hd__a32o_1 _14634_ (.A1(net258),
    .A2(_05623_),
    .A3(_05624_),
    .B1(_05577_),
    .B2(_05578_),
    .X(_08670_));
 sky130_fd_sc_hd__mux2_2 _14635_ (.A0(_04143_),
    .A1(_04145_),
    .S(net305),
    .X(_05625_));
 sky130_fd_sc_hd__nand2_1 _14636_ (.A(net538),
    .B(_05625_),
    .Y(_05626_));
 sky130_fd_sc_hd__a31o_1 _14637_ (.A1(net570),
    .A2(_03010_),
    .A3(_04527_),
    .B1(_03685_),
    .X(_05627_));
 sky130_fd_sc_hd__nand2_1 _14638_ (.A(_05616_),
    .B(_05624_),
    .Y(_05628_));
 sky130_fd_sc_hd__a22oi_1 _14639_ (.A1(net330),
    .A2(net637),
    .B1(net646),
    .B2(net319),
    .Y(_05629_));
 sky130_fd_sc_hd__nand2_4 _14640_ (.A(net319),
    .B(net637),
    .Y(_05631_));
 sky130_fd_sc_hd__and4_2 _14641_ (.A(net319),
    .B(net330),
    .C(net637),
    .D(net646),
    .X(_05632_));
 sky130_fd_sc_hd__nor2_1 _14642_ (.A(_05629_),
    .B(_05632_),
    .Y(_05633_));
 sky130_fd_sc_hd__a21oi_1 _14643_ (.A1(net336),
    .A2(net628),
    .B1(_05633_),
    .Y(_05634_));
 sky130_fd_sc_hd__and3_2 _14644_ (.A(net336),
    .B(net628),
    .C(_05633_),
    .X(_05635_));
 sky130_fd_sc_hd__nor2_1 _14645_ (.A(_05634_),
    .B(_05635_),
    .Y(_05636_));
 sky130_fd_sc_hd__nand2_4 _14646_ (.A(_05590_),
    .B(_05593_),
    .Y(_05637_));
 sky130_fd_sc_hd__o21bai_4 _14647_ (.A1(_05579_),
    .A2(_05583_),
    .B1_N(_05580_),
    .Y(_05638_));
 sky130_fd_sc_hd__and3_2 _14648_ (.A(net343),
    .B(net620),
    .C(_05534_),
    .X(_05639_));
 sky130_fd_sc_hd__xnor2_4 _14649_ (.A(_05638_),
    .B(_05639_),
    .Y(_05640_));
 sky130_fd_sc_hd__inv_2 _14650_ (.A(_05640_),
    .Y(_05642_));
 sky130_fd_sc_hd__xnor2_4 _14651_ (.A(_05637_),
    .B(_05640_),
    .Y(_05643_));
 sky130_fd_sc_hd__nor2_1 _14652_ (.A(_05596_),
    .B(_05600_),
    .Y(_05644_));
 sky130_fd_sc_hd__xnor2_1 _14653_ (.A(_05643_),
    .B(_05644_),
    .Y(_05645_));
 sky130_fd_sc_hd__nand2_1 _14654_ (.A(_05636_),
    .B(_05645_),
    .Y(_05646_));
 sky130_fd_sc_hd__or2_1 _14655_ (.A(_05636_),
    .B(_05645_),
    .X(_05647_));
 sky130_fd_sc_hd__and2_1 _14656_ (.A(_05646_),
    .B(_05647_),
    .X(_05648_));
 sky130_fd_sc_hd__o21ai_2 _14657_ (.A1(_05603_),
    .A2(_05606_),
    .B1(_05648_),
    .Y(_05649_));
 sky130_fd_sc_hd__or3_1 _14658_ (.A(_05603_),
    .B(_05606_),
    .C(_05648_),
    .X(_05650_));
 sky130_fd_sc_hd__and2_4 _14659_ (.A(_05649_),
    .B(_05650_),
    .X(_05651_));
 sky130_fd_sc_hd__nor2_2 _14660_ (.A(_05610_),
    .B(_05613_),
    .Y(_05653_));
 sky130_fd_sc_hd__nand2_1 _14661_ (.A(_05610_),
    .B(_05651_),
    .Y(_05654_));
 sky130_fd_sc_hd__xnor2_4 _14662_ (.A(_05651_),
    .B(_05653_),
    .Y(_05655_));
 sky130_fd_sc_hd__nand2_1 _14663_ (.A(_05628_),
    .B(_05655_),
    .Y(_05656_));
 sky130_fd_sc_hd__or2_1 _14664_ (.A(_05628_),
    .B(_05655_),
    .X(_05657_));
 sky130_fd_sc_hd__a32o_1 _14665_ (.A1(net258),
    .A2(_05656_),
    .A3(_05657_),
    .B1(_05626_),
    .B2(_05627_),
    .X(_08671_));
 sky130_fd_sc_hd__mux2_2 _14666_ (.A0(_04271_),
    .A1(_04273_),
    .S(net305),
    .X(_05658_));
 sky130_fd_sc_hd__nand2_1 _14667_ (.A(net538),
    .B(_05658_),
    .Y(_05659_));
 sky130_fd_sc_hd__a31o_1 _14668_ (.A1(net569),
    .A2(_03186_),
    .A3(_04527_),
    .B1(_03685_),
    .X(_05660_));
 sky130_fd_sc_hd__and2b_1 _14669_ (.A_N(_05616_),
    .B(_05655_),
    .X(_05661_));
 sky130_fd_sc_hd__a31o_1 _14670_ (.A1(_05618_),
    .A2(_05621_),
    .A3(_05655_),
    .B1(_05661_),
    .X(_05663_));
 sky130_fd_sc_hd__a21o_1 _14671_ (.A1(_05613_),
    .A2(_05651_),
    .B1(_05663_),
    .X(_05664_));
 sky130_fd_sc_hd__a31oi_4 _14672_ (.A1(_05618_),
    .A2(_05619_),
    .A3(_05655_),
    .B1(_05664_),
    .Y(_05665_));
 sky130_fd_sc_hd__nand2_8 _14673_ (.A(net330),
    .B(net628),
    .Y(_05666_));
 sky130_fd_sc_hd__or2_2 _14674_ (.A(_05631_),
    .B(_05666_),
    .X(_05667_));
 sky130_fd_sc_hd__xnor2_4 _14675_ (.A(_05631_),
    .B(_05666_),
    .Y(_05668_));
 sky130_fd_sc_hd__nand2_2 _14676_ (.A(net336),
    .B(net620),
    .Y(_05669_));
 sky130_fd_sc_hd__xnor2_1 _14677_ (.A(_05668_),
    .B(_05669_),
    .Y(_05670_));
 sky130_fd_sc_hd__nor2_4 _14678_ (.A(_05632_),
    .B(_05635_),
    .Y(_05671_));
 sky130_fd_sc_hd__nand2b_2 _14679_ (.A_N(_05638_),
    .B(_05534_),
    .Y(_05672_));
 sky130_fd_sc_hd__nand3_4 _14680_ (.A(net343),
    .B(net621),
    .C(_05672_),
    .Y(_05674_));
 sky130_fd_sc_hd__nor2_1 _14681_ (.A(_05671_),
    .B(_05674_),
    .Y(_05675_));
 sky130_fd_sc_hd__xnor2_4 _14682_ (.A(_05671_),
    .B(_05674_),
    .Y(_05676_));
 sky130_fd_sc_hd__and2_1 _14683_ (.A(_05596_),
    .B(_05643_),
    .X(_05677_));
 sky130_fd_sc_hd__inv_2 _14684_ (.A(_05677_),
    .Y(_05678_));
 sky130_fd_sc_hd__a21oi_1 _14685_ (.A1(_05637_),
    .A2(_05642_),
    .B1(_05677_),
    .Y(_05679_));
 sky130_fd_sc_hd__xnor2_1 _14686_ (.A(_05676_),
    .B(_05679_),
    .Y(_05680_));
 sky130_fd_sc_hd__or2_1 _14687_ (.A(_05670_),
    .B(_05680_),
    .X(_05681_));
 sky130_fd_sc_hd__nand2_1 _14688_ (.A(_05670_),
    .B(_05680_),
    .Y(_05682_));
 sky130_fd_sc_hd__nand2_1 _14689_ (.A(_05681_),
    .B(_05682_),
    .Y(_05683_));
 sky130_fd_sc_hd__nor2_1 _14690_ (.A(_05646_),
    .B(_05683_),
    .Y(_05685_));
 sky130_fd_sc_hd__and2_1 _14691_ (.A(_05646_),
    .B(_05683_),
    .X(_05686_));
 sky130_fd_sc_hd__nor2_1 _14692_ (.A(_05685_),
    .B(_05686_),
    .Y(_05687_));
 sky130_fd_sc_hd__and3_1 _14693_ (.A(_05600_),
    .B(_05643_),
    .C(_05687_),
    .X(_05688_));
 sky130_fd_sc_hd__a21oi_1 _14694_ (.A1(_05600_),
    .A2(_05643_),
    .B1(_05687_),
    .Y(_05689_));
 sky130_fd_sc_hd__or2_2 _14695_ (.A(_05688_),
    .B(_05689_),
    .X(_05690_));
 sky130_fd_sc_hd__nor2_1 _14696_ (.A(_05649_),
    .B(_05690_),
    .Y(_05691_));
 sky130_fd_sc_hd__nor2_1 _14697_ (.A(_05654_),
    .B(_05690_),
    .Y(_05692_));
 sky130_fd_sc_hd__nand2_1 _14698_ (.A(_05649_),
    .B(_05654_),
    .Y(_05693_));
 sky130_fd_sc_hd__xor2_2 _14699_ (.A(_05690_),
    .B(_05693_),
    .X(_05694_));
 sky130_fd_sc_hd__nand2_1 _14700_ (.A(_05665_),
    .B(_05694_),
    .Y(_05696_));
 sky130_fd_sc_hd__nor2_1 _14701_ (.A(_05665_),
    .B(_05694_),
    .Y(_05697_));
 sky130_fd_sc_hd__inv_2 _14702_ (.A(_05697_),
    .Y(_05698_));
 sky130_fd_sc_hd__a32o_1 _14703_ (.A1(net259),
    .A2(_05696_),
    .A3(_05698_),
    .B1(_05659_),
    .B2(_05660_),
    .X(_08672_));
 sky130_fd_sc_hd__mux2_2 _14704_ (.A0(_04408_),
    .A1(_04410_),
    .S(net306),
    .X(_05699_));
 sky130_fd_sc_hd__nand2_1 _14705_ (.A(net539),
    .B(_05699_),
    .Y(_05700_));
 sky130_fd_sc_hd__a31o_1 _14706_ (.A1(net570),
    .A2(_03353_),
    .A3(_04527_),
    .B1(_03685_),
    .X(_05701_));
 sky130_fd_sc_hd__a22o_1 _14707_ (.A1(net329),
    .A2(net620),
    .B1(net628),
    .B2(net320),
    .X(_05702_));
 sky130_fd_sc_hd__nand4_1 _14708_ (.A(net320),
    .B(net329),
    .C(net620),
    .D(net628),
    .Y(_05703_));
 sky130_fd_sc_hd__o21ai_4 _14709_ (.A1(_05668_),
    .A2(_05669_),
    .B1(_05667_),
    .Y(_05704_));
 sky130_fd_sc_hd__and3b_1 _14710_ (.A_N(_05676_),
    .B(_05642_),
    .C(_05637_),
    .X(_05706_));
 sky130_fd_sc_hd__nor2_1 _14711_ (.A(_05675_),
    .B(_05706_),
    .Y(_05707_));
 sky130_fd_sc_hd__xnor2_2 _14712_ (.A(_05704_),
    .B(_05707_),
    .Y(_05708_));
 sky130_fd_sc_hd__nand3_1 _14713_ (.A(_05702_),
    .B(_05703_),
    .C(_05708_),
    .Y(_05709_));
 sky130_fd_sc_hd__a21o_1 _14714_ (.A1(_05702_),
    .A2(_05703_),
    .B1(_05708_),
    .X(_05710_));
 sky130_fd_sc_hd__nand2_1 _14715_ (.A(_05709_),
    .B(_05710_),
    .Y(_05711_));
 sky130_fd_sc_hd__or2_1 _14716_ (.A(_05681_),
    .B(_05711_),
    .X(_05712_));
 sky130_fd_sc_hd__nand2_1 _14717_ (.A(_05681_),
    .B(_05711_),
    .Y(_05713_));
 sky130_fd_sc_hd__nand2_1 _14718_ (.A(_05712_),
    .B(_05713_),
    .Y(_05714_));
 sky130_fd_sc_hd__or3_1 _14719_ (.A(_05676_),
    .B(_05678_),
    .C(_05714_),
    .X(_05715_));
 sky130_fd_sc_hd__o21ai_1 _14720_ (.A1(_05676_),
    .A2(_05678_),
    .B1(_05714_),
    .Y(_05717_));
 sky130_fd_sc_hd__and2_1 _14721_ (.A(_05715_),
    .B(_05717_),
    .X(_05718_));
 sky130_fd_sc_hd__o21ai_2 _14722_ (.A1(_05685_),
    .A2(_05688_),
    .B1(_05718_),
    .Y(_05719_));
 sky130_fd_sc_hd__or3_1 _14723_ (.A(_05685_),
    .B(_05688_),
    .C(_05718_),
    .X(_05720_));
 sky130_fd_sc_hd__and2_1 _14724_ (.A(_05719_),
    .B(_05720_),
    .X(_05721_));
 sky130_fd_sc_hd__inv_2 _14725_ (.A(_05721_),
    .Y(_05722_));
 sky130_fd_sc_hd__and3_1 _14726_ (.A(_05691_),
    .B(_05719_),
    .C(_05720_),
    .X(_05723_));
 sky130_fd_sc_hd__or2_1 _14727_ (.A(_05691_),
    .B(_05721_),
    .X(_05724_));
 sky130_fd_sc_hd__nand2b_1 _14728_ (.A_N(_05723_),
    .B(_05724_),
    .Y(_05725_));
 sky130_fd_sc_hd__nor2_1 _14729_ (.A(_05692_),
    .B(_05697_),
    .Y(_05726_));
 sky130_fd_sc_hd__nand2_1 _14730_ (.A(_05725_),
    .B(_05726_),
    .Y(_05728_));
 sky130_fd_sc_hd__or2_1 _14731_ (.A(_05725_),
    .B(_05726_),
    .X(_05729_));
 sky130_fd_sc_hd__a32o_1 _14732_ (.A1(net258),
    .A2(_05728_),
    .A3(_05729_),
    .B1(_05700_),
    .B2(_05701_),
    .X(_08673_));
 sky130_fd_sc_hd__mux2_1 _14733_ (.A0(_04525_),
    .A1(_04529_),
    .S(net308),
    .X(_05730_));
 sky130_fd_sc_hd__nand2_1 _14734_ (.A(net538),
    .B(_05730_),
    .Y(_05731_));
 sky130_fd_sc_hd__a31o_1 _14735_ (.A1(net570),
    .A2(_03518_),
    .A3(_04527_),
    .B1(_03685_),
    .X(_05732_));
 sky130_fd_sc_hd__nand2_1 _14736_ (.A(_05675_),
    .B(_05704_),
    .Y(_05733_));
 sky130_fd_sc_hd__or2_1 _14737_ (.A(_05666_),
    .B(_05733_),
    .X(_05734_));
 sky130_fd_sc_hd__nand2_2 _14738_ (.A(net319),
    .B(net620),
    .Y(_05735_));
 sky130_fd_sc_hd__nand2_1 _14739_ (.A(_05666_),
    .B(_05733_),
    .Y(_05736_));
 sky130_fd_sc_hd__o21a_1 _14740_ (.A1(_05735_),
    .A2(_05736_),
    .B1(_05734_),
    .X(_05738_));
 sky130_fd_sc_hd__or2_1 _14741_ (.A(_05709_),
    .B(_05738_),
    .X(_05739_));
 sky130_fd_sc_hd__nand2_1 _14742_ (.A(_05709_),
    .B(_05738_),
    .Y(_05740_));
 sky130_fd_sc_hd__nand2_1 _14743_ (.A(_05739_),
    .B(_05740_),
    .Y(_05741_));
 sky130_fd_sc_hd__nand2_1 _14744_ (.A(_05704_),
    .B(_05706_),
    .Y(_05742_));
 sky130_fd_sc_hd__xnor2_1 _14745_ (.A(_05741_),
    .B(_05742_),
    .Y(_05743_));
 sky130_fd_sc_hd__a21oi_1 _14746_ (.A1(_05712_),
    .A2(_05715_),
    .B1(_05743_),
    .Y(_05744_));
 sky130_fd_sc_hd__and3_1 _14747_ (.A(_05712_),
    .B(_05715_),
    .C(_05743_),
    .X(_05745_));
 sky130_fd_sc_hd__or2_1 _14748_ (.A(_05744_),
    .B(_05745_),
    .X(_05746_));
 sky130_fd_sc_hd__or2_1 _14749_ (.A(_05719_),
    .B(_05746_),
    .X(_05747_));
 sky130_fd_sc_hd__nand2_1 _14750_ (.A(_05719_),
    .B(_05746_),
    .Y(_05749_));
 sky130_fd_sc_hd__nand2_1 _14751_ (.A(_05747_),
    .B(_05749_),
    .Y(_05750_));
 sky130_fd_sc_hd__o21ai_1 _14752_ (.A1(_05692_),
    .A2(_05723_),
    .B1(_05724_),
    .Y(_05751_));
 sky130_fd_sc_hd__o31a_1 _14753_ (.A1(_05665_),
    .A2(_05694_),
    .A3(_05722_),
    .B1(_05751_),
    .X(_05752_));
 sky130_fd_sc_hd__nand2_1 _14754_ (.A(_05750_),
    .B(_05752_),
    .Y(_05753_));
 sky130_fd_sc_hd__or2_1 _14755_ (.A(_05750_),
    .B(_05752_),
    .X(_05754_));
 sky130_fd_sc_hd__a32o_1 _14756_ (.A1(net259),
    .A2(_05753_),
    .A3(_05754_),
    .B1(_05731_),
    .B2(_05732_),
    .X(_08674_));
 sky130_fd_sc_hd__mux2_1 _14757_ (.A0(_04753_),
    .A1(_04755_),
    .S(net305),
    .X(_05755_));
 sky130_fd_sc_hd__nor2_1 _14758_ (.A(_03686_),
    .B(_05755_),
    .Y(_05756_));
 sky130_fd_sc_hd__o21a_1 _14759_ (.A1(_05750_),
    .A2(_05752_),
    .B1(_05747_),
    .X(_05757_));
 sky130_fd_sc_hd__o21ai_1 _14760_ (.A1(_05741_),
    .A2(_05742_),
    .B1(_05739_),
    .Y(_05759_));
 sky130_fd_sc_hd__a311o_1 _14761_ (.A1(net320),
    .A2(net621),
    .A3(_05736_),
    .B1(_05744_),
    .C1(_05759_),
    .X(_05760_));
 sky130_fd_sc_hd__xnor2_1 _14762_ (.A(_05757_),
    .B(_05760_),
    .Y(_05761_));
 sky130_fd_sc_hd__mux2_1 _14763_ (.A0(_05756_),
    .A1(_05761_),
    .S(net259),
    .X(_08676_));
 sky130_fd_sc_hd__nor2_1 _14764_ (.A(net343),
    .B(net646),
    .Y(_05762_));
 sky130_fd_sc_hd__or2_1 _14765_ (.A(net343),
    .B(net646),
    .X(_05763_));
 sky130_fd_sc_hd__or2_1 _14766_ (.A(net354),
    .B(net658),
    .X(_05764_));
 sky130_fd_sc_hd__nor2_1 _14767_ (.A(net361),
    .B(net666),
    .Y(_05765_));
 sky130_fd_sc_hd__or2_1 _14768_ (.A(net361),
    .B(net666),
    .X(_05766_));
 sky130_fd_sc_hd__or2_4 _14769_ (.A(net370),
    .B(net674),
    .X(_05767_));
 sky130_fd_sc_hd__or2_1 _14770_ (.A(net379),
    .B(net678),
    .X(_05769_));
 sky130_fd_sc_hd__or2_1 _14771_ (.A(net386),
    .B(net688),
    .X(_05770_));
 sky130_fd_sc_hd__or2_1 _14772_ (.A(net395),
    .B(net697),
    .X(_05771_));
 sky130_fd_sc_hd__or2_2 _14773_ (.A(net402),
    .B(net709),
    .X(_05772_));
 sky130_fd_sc_hd__or2_1 _14774_ (.A(net410),
    .B(net717),
    .X(_05773_));
 sky130_fd_sc_hd__or2_2 _14775_ (.A(net417),
    .B(net727),
    .X(_05774_));
 sky130_fd_sc_hd__or2_1 _14776_ (.A(net426),
    .B(net735),
    .X(_05775_));
 sky130_fd_sc_hd__or2_2 _14777_ (.A(net434),
    .B(net744),
    .X(_05776_));
 sky130_fd_sc_hd__or2_2 _14778_ (.A(net444),
    .B(net753),
    .X(_05777_));
 sky130_fd_sc_hd__or2_2 _14779_ (.A(net451),
    .B(net764),
    .X(_05778_));
 sky130_fd_sc_hd__or2_2 _14780_ (.A(net461),
    .B(net774),
    .X(_05780_));
 sky130_fd_sc_hd__or2_2 _14781_ (.A(net471),
    .B(net786),
    .X(_05781_));
 sky130_fd_sc_hd__or2_1 _14782_ (.A(net478),
    .B(net798),
    .X(_05782_));
 sky130_fd_sc_hd__or2_2 _14783_ (.A(net490),
    .B(net807),
    .X(_05783_));
 sky130_fd_sc_hd__or2_1 _14784_ (.A(net499),
    .B(net816),
    .X(_05784_));
 sky130_fd_sc_hd__or2_2 _14785_ (.A(net507),
    .B(net827),
    .X(_05785_));
 sky130_fd_sc_hd__or2_1 _14786_ (.A(net514),
    .B(net836),
    .X(_05786_));
 sky130_fd_sc_hd__nor2_2 _14787_ (.A(net523),
    .B(net847),
    .Y(_05787_));
 sky130_fd_sc_hd__nor2_1 _14788_ (.A(net532),
    .B(net857),
    .Y(_05788_));
 sky130_fd_sc_hd__nor2_1 _14789_ (.A(net545),
    .B(net865),
    .Y(_05789_));
 sky130_fd_sc_hd__nor2_1 _14790_ (.A(net560),
    .B(net876),
    .Y(_05791_));
 sky130_fd_sc_hd__or2_2 _14791_ (.A(net578),
    .B(net886),
    .X(_05792_));
 sky130_fd_sc_hd__or2_2 _14792_ (.A(net590),
    .B(net898),
    .X(_05793_));
 sky130_fd_sc_hd__nor2_1 _14793_ (.A(net603),
    .B(net906),
    .Y(_05794_));
 sky130_fd_sc_hd__or2_2 _14794_ (.A(net603),
    .B(net905),
    .X(_05795_));
 sky130_fd_sc_hd__a22o_1 _14795_ (.A1(net603),
    .A2(net906),
    .B1(net914),
    .B2(net615),
    .X(_05796_));
 sky130_fd_sc_hd__and4_1 _14796_ (.A(_02387_),
    .B(_05793_),
    .C(_05795_),
    .D(_05796_),
    .X(_05797_));
 sky130_fd_sc_hd__a31o_2 _14797_ (.A1(_05793_),
    .A2(_05795_),
    .A3(_05796_),
    .B1(_02386_),
    .X(_05798_));
 sky130_fd_sc_hd__a21oi_2 _14798_ (.A1(_05792_),
    .A2(_05798_),
    .B1(_02264_),
    .Y(_05799_));
 sky130_fd_sc_hd__o21ba_1 _14799_ (.A1(_05791_),
    .A2(_05799_),
    .B1_N(_02116_),
    .X(_05800_));
 sky130_fd_sc_hd__o21ba_1 _14800_ (.A1(_05789_),
    .A2(_05800_),
    .B1_N(_02060_),
    .X(_05802_));
 sky130_fd_sc_hd__or3_1 _14801_ (.A(_01662_),
    .B(_05788_),
    .C(_05802_),
    .X(_05803_));
 sky130_fd_sc_hd__o21a_1 _14802_ (.A1(_05788_),
    .A2(_05802_),
    .B1(_01663_),
    .X(_05804_));
 sky130_fd_sc_hd__nor2_1 _14803_ (.A(_05787_),
    .B(_05804_),
    .Y(_05805_));
 sky130_fd_sc_hd__o21ai_1 _14804_ (.A1(_05787_),
    .A2(_05804_),
    .B1(_01594_),
    .Y(_05806_));
 sky130_fd_sc_hd__and3_1 _14805_ (.A(_01716_),
    .B(_05786_),
    .C(_05806_),
    .X(_05807_));
 sky130_fd_sc_hd__or2_2 _14806_ (.A(_01715_),
    .B(_05807_),
    .X(_05808_));
 sky130_fd_sc_hd__a21bo_2 _14807_ (.A1(_05785_),
    .A2(_05808_),
    .B1_N(_01414_),
    .X(_05809_));
 sky130_fd_sc_hd__a21o_1 _14808_ (.A1(_05784_),
    .A2(_05809_),
    .B1(_01064_),
    .X(_05810_));
 sky130_fd_sc_hd__a21o_2 _14809_ (.A1(_05783_),
    .A2(_05810_),
    .B1(_00936_),
    .X(_05811_));
 sky130_fd_sc_hd__a21o_1 _14810_ (.A1(_05782_),
    .A2(_05811_),
    .B1(_00653_),
    .X(_05813_));
 sky130_fd_sc_hd__a21o_1 _14811_ (.A1(_05781_),
    .A2(_05813_),
    .B1(_00219_),
    .X(_05814_));
 sky130_fd_sc_hd__a21bo_1 _14812_ (.A1(_05780_),
    .A2(_05814_),
    .B1_N(_08626_),
    .X(_05815_));
 sky130_fd_sc_hd__a21bo_1 _14813_ (.A1(_05778_),
    .A2(_05815_),
    .B1_N(_05001_),
    .X(_05816_));
 sky130_fd_sc_hd__a21o_1 _14814_ (.A1(_05777_),
    .A2(_05816_),
    .B1(_03637_),
    .X(_05817_));
 sky130_fd_sc_hd__a21bo_1 _14815_ (.A1(_05776_),
    .A2(_05817_),
    .B1_N(_03659_),
    .X(_05818_));
 sky130_fd_sc_hd__a21o_1 _14816_ (.A1(_05775_),
    .A2(_05818_),
    .B1(_03025_),
    .X(_05819_));
 sky130_fd_sc_hd__a21bo_1 _14817_ (.A1(_05774_),
    .A2(_05819_),
    .B1_N(_03363_),
    .X(_05820_));
 sky130_fd_sc_hd__a21o_1 _14818_ (.A1(_05773_),
    .A2(_05820_),
    .B1(_03365_),
    .X(_05821_));
 sky130_fd_sc_hd__a21bo_1 _14819_ (.A1(_05772_),
    .A2(_05821_),
    .B1_N(_04070_),
    .X(_05822_));
 sky130_fd_sc_hd__a21o_1 _14820_ (.A1(_05771_),
    .A2(_05822_),
    .B1(_04334_),
    .X(_05824_));
 sky130_fd_sc_hd__a21bo_1 _14821_ (.A1(_05770_),
    .A2(_05824_),
    .B1_N(_04597_),
    .X(_05825_));
 sky130_fd_sc_hd__a21bo_2 _14822_ (.A1(_05769_),
    .A2(_05825_),
    .B1_N(_04820_),
    .X(_05826_));
 sky130_fd_sc_hd__a21oi_4 _14823_ (.A1(_05767_),
    .A2(_05826_),
    .B1(_04928_),
    .Y(_05827_));
 sky130_fd_sc_hd__o21ai_2 _14824_ (.A1(_05765_),
    .A2(_05827_),
    .B1(_05182_),
    .Y(_05828_));
 sky130_fd_sc_hd__nand2_1 _14825_ (.A(_05764_),
    .B(_05828_),
    .Y(_05829_));
 sky130_fd_sc_hd__a211o_2 _14826_ (.A1(_05334_),
    .A2(_05829_),
    .B1(_05762_),
    .C1(_05408_),
    .X(_05830_));
 sky130_fd_sc_hd__nor2_2 _14827_ (.A(net336),
    .B(net638),
    .Y(_05831_));
 sky130_fd_sc_hd__a211oi_4 _14828_ (.A1(_05407_),
    .A2(_05830_),
    .B1(_05831_),
    .C1(_05582_),
    .Y(_05832_));
 sky130_fd_sc_hd__or2_4 _14829_ (.A(net329),
    .B(net628),
    .X(_05833_));
 sky130_fd_sc_hd__o211ai_4 _14830_ (.A1(_05582_),
    .A2(_05832_),
    .B1(_05833_),
    .C1(_05666_),
    .Y(_05835_));
 sky130_fd_sc_hd__nand3_1 _14831_ (.A(_05666_),
    .B(_05735_),
    .C(_05835_),
    .Y(_05836_));
 sky130_fd_sc_hd__or2_1 _14832_ (.A(net319),
    .B(net620),
    .X(_05837_));
 sky130_fd_sc_hd__or2_4 _14833_ (.A(net316),
    .B(net315),
    .X(_05838_));
 sky130_fd_sc_hd__nand2b_4 _14834_ (.A_N(net315),
    .B(net316),
    .Y(_05839_));
 sky130_fd_sc_hd__and3_4 _14835_ (.A(net277),
    .B(_03367_),
    .C(_05838_),
    .X(_05840_));
 sky130_fd_sc_hd__nand3_2 _14836_ (.A(net277),
    .B(_03367_),
    .C(_05838_),
    .Y(_05841_));
 sky130_fd_sc_hd__nor2_1 _14837_ (.A(_02576_),
    .B(net255),
    .Y(_05842_));
 sky130_fd_sc_hd__o21a_2 _14838_ (.A1(_00621_),
    .A2(_02574_),
    .B1(_05842_),
    .X(_05843_));
 sky130_fd_sc_hd__nor2_1 _14839_ (.A(net553),
    .B(_04762_),
    .Y(_05844_));
 sky130_fd_sc_hd__nor2_1 _14840_ (.A(net308),
    .B(_04759_),
    .Y(_05846_));
 sky130_fd_sc_hd__nor2_1 _14841_ (.A(net207),
    .B(_04758_),
    .Y(_05847_));
 sky130_fd_sc_hd__o32a_1 _14842_ (.A1(net537),
    .A2(_05844_),
    .A3(_05846_),
    .B1(_05847_),
    .B2(_02643_),
    .X(_05848_));
 sky130_fd_sc_hd__nor2_4 _14843_ (.A(_03388_),
    .B(_05839_),
    .Y(_05849_));
 sky130_fd_sc_hd__or2_4 _14844_ (.A(_03388_),
    .B(_05839_),
    .X(_05850_));
 sky130_fd_sc_hd__nand2_1 _14845_ (.A(net905),
    .B(net914),
    .Y(_05851_));
 sky130_fd_sc_hd__nor2_2 _14846_ (.A(_03280_),
    .B(_05851_),
    .Y(_05852_));
 sky130_fd_sc_hd__and2_1 _14847_ (.A(net886),
    .B(_05852_),
    .X(_05853_));
 sky130_fd_sc_hd__and3_1 _14848_ (.A(net868),
    .B(net875),
    .C(_05853_),
    .X(_05854_));
 sky130_fd_sc_hd__and2_1 _14849_ (.A(net855),
    .B(_05854_),
    .X(_05855_));
 sky130_fd_sc_hd__and3_1 _14850_ (.A(net845),
    .B(net855),
    .C(_05854_),
    .X(_05857_));
 sky130_fd_sc_hd__and2_1 _14851_ (.A(net838),
    .B(_05857_),
    .X(_05858_));
 sky130_fd_sc_hd__and3_1 _14852_ (.A(net827),
    .B(net838),
    .C(_05857_),
    .X(_05859_));
 sky130_fd_sc_hd__and3_2 _14853_ (.A(net816),
    .B(net829),
    .C(_05858_),
    .X(_05860_));
 sky130_fd_sc_hd__and2_1 _14854_ (.A(net807),
    .B(_05860_),
    .X(_05861_));
 sky130_fd_sc_hd__and3_1 _14855_ (.A(net796),
    .B(net807),
    .C(_05860_),
    .X(_05862_));
 sky130_fd_sc_hd__and3_1 _14856_ (.A(net786),
    .B(net796),
    .C(_05861_),
    .X(_05863_));
 sky130_fd_sc_hd__and2_1 _14857_ (.A(net775),
    .B(_05863_),
    .X(_05864_));
 sky130_fd_sc_hd__and3_2 _14858_ (.A(net764),
    .B(net775),
    .C(_05863_),
    .X(_05865_));
 sky130_fd_sc_hd__and3_1 _14859_ (.A(net744),
    .B(net753),
    .C(_05865_),
    .X(_05866_));
 sky130_fd_sc_hd__and2_2 _14860_ (.A(net735),
    .B(_05866_),
    .X(_05868_));
 sky130_fd_sc_hd__and3_1 _14861_ (.A(net717),
    .B(net727),
    .C(_05868_),
    .X(_05869_));
 sky130_fd_sc_hd__and2_2 _14862_ (.A(net709),
    .B(_05869_),
    .X(_05870_));
 sky130_fd_sc_hd__and3_1 _14863_ (.A(net688),
    .B(net697),
    .C(_05870_),
    .X(_05871_));
 sky130_fd_sc_hd__and2_2 _14864_ (.A(net678),
    .B(_05871_),
    .X(_05872_));
 sky130_fd_sc_hd__and3_1 _14865_ (.A(net666),
    .B(net674),
    .C(_05872_),
    .X(_05873_));
 sky130_fd_sc_hd__and2_2 _14866_ (.A(net658),
    .B(_05873_),
    .X(_05874_));
 sky130_fd_sc_hd__and3_1 _14867_ (.A(net637),
    .B(net646),
    .C(_05874_),
    .X(_05875_));
 sky130_fd_sc_hd__and2_1 _14868_ (.A(net628),
    .B(_05875_),
    .X(_05876_));
 sky130_fd_sc_hd__a311o_1 _14869_ (.A1(net618),
    .A2(_05849_),
    .A3(_05876_),
    .B1(_05843_),
    .C1(_05848_),
    .X(_05877_));
 sky130_fd_sc_hd__a31o_1 _14870_ (.A1(_05836_),
    .A2(_05837_),
    .A3(_05840_),
    .B1(_05877_),
    .X(_08716_));
 sky130_fd_sc_hd__nor2_1 _14871_ (.A(_03452_),
    .B(_05838_),
    .Y(_05879_));
 sky130_fd_sc_hd__or2_4 _14872_ (.A(_03452_),
    .B(_05838_),
    .X(_05880_));
 sky130_fd_sc_hd__or3b_2 _14873_ (.A(net451),
    .B(net461),
    .C_N(net310),
    .X(_05881_));
 sky130_fd_sc_hd__or3_2 _14874_ (.A(net500),
    .B(_02587_),
    .C(_05881_),
    .X(_05882_));
 sky130_fd_sc_hd__or3_1 _14875_ (.A(_02587_),
    .B(_02588_),
    .C(_05881_),
    .X(_05883_));
 sky130_fd_sc_hd__or4_1 _14876_ (.A(net515),
    .B(_02587_),
    .C(_02588_),
    .D(_05881_),
    .X(_05884_));
 sky130_fd_sc_hd__o21bai_4 _14877_ (.A1(\sel_op[3] ),
    .A2(net311),
    .B1_N(net310),
    .Y(_05885_));
 sky130_fd_sc_hd__a21o_1 _14878_ (.A1(net311),
    .A2(_02583_),
    .B1(_05885_),
    .X(_05886_));
 sky130_fd_sc_hd__nand2b_1 _14879_ (.A_N(net311),
    .B(\sel_op[3] ),
    .Y(_05887_));
 sky130_fd_sc_hd__a21o_1 _14880_ (.A1(net311),
    .A2(_02586_),
    .B1(_05885_),
    .X(_05889_));
 sky130_fd_sc_hd__a21o_4 _14881_ (.A1(_05884_),
    .A2(_05889_),
    .B1(net312),
    .X(_05890_));
 sky130_fd_sc_hd__or3_2 _14882_ (.A(net490),
    .B(_03335_),
    .C(_02586_),
    .X(_05891_));
 sky130_fd_sc_hd__or3b_1 _14883_ (.A(net500),
    .B(net507),
    .C_N(net312),
    .X(_05892_));
 sky130_fd_sc_hd__or3_4 _14884_ (.A(_02583_),
    .B(_02587_),
    .C(_05892_),
    .X(_05893_));
 sky130_fd_sc_hd__or4_2 _14885_ (.A(net515),
    .B(_02583_),
    .C(_02587_),
    .D(_05892_),
    .X(_05894_));
 sky130_fd_sc_hd__or4_2 _14886_ (.A(net523),
    .B(net533),
    .C(net547),
    .D(_05894_),
    .X(_05895_));
 sky130_fd_sc_hd__nor2_2 _14887_ (.A(_02582_),
    .B(_05893_),
    .Y(_05896_));
 sky130_fd_sc_hd__or4_2 _14888_ (.A(_02582_),
    .B(_02583_),
    .C(_02587_),
    .D(_05892_),
    .X(_05897_));
 sky130_fd_sc_hd__or4_4 _14889_ (.A(net533),
    .B(net547),
    .C(net562),
    .D(_05897_),
    .X(_05898_));
 sky130_fd_sc_hd__a21oi_1 _14890_ (.A1(_05890_),
    .A2(_05898_),
    .B1(net286),
    .Y(_05900_));
 sky130_fd_sc_hd__a21o_4 _14891_ (.A1(_05890_),
    .A2(_05898_),
    .B1(net286),
    .X(_05901_));
 sky130_fd_sc_hd__or3_4 _14892_ (.A(net763),
    .B(net774),
    .C(net785),
    .X(_05902_));
 sky130_fd_sc_hd__or2_1 _14893_ (.A(net796),
    .B(net808),
    .X(_05903_));
 sky130_fd_sc_hd__or3_4 _14894_ (.A(net796),
    .B(net807),
    .C(net818),
    .X(_05904_));
 sky130_fd_sc_hd__or2_1 _14895_ (.A(net828),
    .B(net837),
    .X(_05905_));
 sky130_fd_sc_hd__or3b_1 _14896_ (.A(net828),
    .B(net848),
    .C_N(net313),
    .X(_05906_));
 sky130_fd_sc_hd__or4_4 _14897_ (.A(net837),
    .B(_05902_),
    .C(_05904_),
    .D(_05906_),
    .X(_05907_));
 sky130_fd_sc_hd__inv_2 _14898_ (.A(_05907_),
    .Y(_05908_));
 sky130_fd_sc_hd__or3_4 _14899_ (.A(net858),
    .B(net867),
    .C(_05907_),
    .X(_05909_));
 sky130_fd_sc_hd__o21a_1 _14900_ (.A1(net763),
    .A2(net774),
    .B1(net311),
    .X(_05911_));
 sky130_fd_sc_hd__or2_1 _14901_ (.A(net785),
    .B(net797),
    .X(_05912_));
 sky130_fd_sc_hd__or4b_2 _14902_ (.A(net763),
    .B(net774),
    .C(net785),
    .D_N(net310),
    .X(_05913_));
 sky130_fd_sc_hd__a2111o_1 _14903_ (.A1(_05887_),
    .A2(_05912_),
    .B1(_05911_),
    .C1(net312),
    .D1(_05885_),
    .X(_05914_));
 sky130_fd_sc_hd__nand2b_1 _14904_ (.A_N(net313),
    .B(net310),
    .Y(_05915_));
 sky130_fd_sc_hd__or4_1 _14905_ (.A(_05902_),
    .B(_05904_),
    .C(_05905_),
    .D(_05915_),
    .X(_05916_));
 sky130_fd_sc_hd__or3_1 _14906_ (.A(net858),
    .B(net867),
    .C(net878),
    .X(_05917_));
 sky130_fd_sc_hd__o211a_4 _14907_ (.A1(_05907_),
    .A2(_05917_),
    .B1(_05916_),
    .C1(_05914_),
    .X(_05918_));
 sky130_fd_sc_hd__nor2_4 _14908_ (.A(_03302_),
    .B(_05918_),
    .Y(_05919_));
 sky130_fd_sc_hd__or2_4 _14909_ (.A(_03302_),
    .B(_05918_),
    .X(_05920_));
 sky130_fd_sc_hd__and3_1 _14910_ (.A(net280),
    .B(net154),
    .C(net153),
    .X(_05922_));
 sky130_fd_sc_hd__and2b_2 _14911_ (.A_N(net527),
    .B(net213),
    .X(_05923_));
 sky130_fd_sc_hd__nand2b_1 _14912_ (.A_N(net527),
    .B(net214),
    .Y(_05924_));
 sky130_fd_sc_hd__a21oi_1 _14913_ (.A1(net284),
    .A2(net771),
    .B1(_01580_),
    .Y(_05925_));
 sky130_fd_sc_hd__mux2_1 _14914_ (.A0(net793),
    .A1(net783),
    .S(net609),
    .X(_05926_));
 sky130_fd_sc_hd__nor2_1 _14915_ (.A(net600),
    .B(_05926_),
    .Y(_05927_));
 sky130_fd_sc_hd__a211o_1 _14916_ (.A1(net601),
    .A2(_05925_),
    .B1(_05927_),
    .C1(net150),
    .X(_05928_));
 sky130_fd_sc_hd__mux4_1 _14917_ (.A0(net838),
    .A1(net829),
    .A2(net819),
    .A3(net807),
    .S0(net610),
    .S1(net601),
    .X(_05929_));
 sky130_fd_sc_hd__nand2_1 _14918_ (.A(net151),
    .B(_05929_),
    .Y(_05930_));
 sky130_fd_sc_hd__mux2_1 _14919_ (.A0(_05928_),
    .A1(_05930_),
    .S(net299),
    .X(_05931_));
 sky130_fd_sc_hd__mux4_1 _14920_ (.A0(net912),
    .A1(net902),
    .A2(net898),
    .A3(net886),
    .S0(net609),
    .S1(net601),
    .X(_05933_));
 sky130_fd_sc_hd__mux4_1 _14921_ (.A0(net875),
    .A1(net868),
    .A2(net855),
    .A3(net845),
    .S0(net610),
    .S1(net601),
    .X(_05934_));
 sky130_fd_sc_hd__mux2_1 _14922_ (.A0(_05933_),
    .A1(_05934_),
    .S(net592),
    .X(_05935_));
 sky130_fd_sc_hd__a21oi_1 _14923_ (.A1(net151),
    .A2(_05935_),
    .B1(net576),
    .Y(_05936_));
 sky130_fd_sc_hd__or3_4 _14924_ (.A(net544),
    .B(_03388_),
    .C(_02577_),
    .X(_05937_));
 sky130_fd_sc_hd__nor2_1 _14925_ (.A(net559),
    .B(_05937_),
    .Y(_05938_));
 sky130_fd_sc_hd__or2_2 _14926_ (.A(net559),
    .B(_05937_),
    .X(_05939_));
 sky130_fd_sc_hd__a211o_2 _14927_ (.A1(net576),
    .A2(_05931_),
    .B1(_05936_),
    .C1(net202),
    .X(_05940_));
 sky130_fd_sc_hd__nor2_1 _14928_ (.A(_03388_),
    .B(_05838_),
    .Y(_05941_));
 sky130_fd_sc_hd__or2_4 _14929_ (.A(_03388_),
    .B(_05838_),
    .X(_05942_));
 sky130_fd_sc_hd__nor3b_2 _14930_ (.A(net316),
    .B(net315),
    .C_N(_03367_),
    .Y(_05944_));
 sky130_fd_sc_hd__or3b_4 _14931_ (.A(net316),
    .B(net315),
    .C_N(_03367_),
    .X(_05945_));
 sky130_fd_sc_hd__a21oi_1 _14932_ (.A1(net255),
    .A2(net235),
    .B1(net285),
    .Y(_05946_));
 sky130_fd_sc_hd__nor2_1 _14933_ (.A(_03420_),
    .B(_05838_),
    .Y(_05947_));
 sky130_fd_sc_hd__a2111o_1 _14934_ (.A1(net285),
    .A2(net254),
    .B1(_05946_),
    .C1(net234),
    .D1(_03302_),
    .X(_05948_));
 sky130_fd_sc_hd__o31a_1 _14935_ (.A1(net912),
    .A2(net254),
    .A3(_05849_),
    .B1(_05948_),
    .X(_05949_));
 sky130_fd_sc_hd__o32a_1 _14936_ (.A1(net611),
    .A2(net912),
    .A3(_05849_),
    .B1(net240),
    .B2(_05949_),
    .X(_05950_));
 sky130_fd_sc_hd__nor2_4 _14937_ (.A(\op_code[0] ),
    .B(_05839_),
    .Y(_05951_));
 sky130_fd_sc_hd__or2_4 _14938_ (.A(\op_code[0] ),
    .B(_05839_),
    .X(_05952_));
 sky130_fd_sc_hd__and4bb_1 _14939_ (.A_N(\op_code[0] ),
    .B_N(\op_code[3] ),
    .C(net316),
    .D(\op_code[1] ),
    .X(_05953_));
 sky130_fd_sc_hd__or4bb_4 _14940_ (.A(\op_code[0] ),
    .B(net315),
    .C_N(net316),
    .D_N(\op_code[1] ),
    .X(_05955_));
 sky130_fd_sc_hd__a21o_1 _14941_ (.A1(net285),
    .A2(net272),
    .B1(net912),
    .X(_05956_));
 sky130_fd_sc_hd__or3_1 _14942_ (.A(net611),
    .B(_03302_),
    .C(net269),
    .X(_05957_));
 sky130_fd_sc_hd__a21oi_1 _14943_ (.A1(_05956_),
    .A2(_05957_),
    .B1(net228),
    .Y(_05958_));
 sky130_fd_sc_hd__nor3_1 _14944_ (.A(net244),
    .B(_05950_),
    .C(_05958_),
    .Y(_05959_));
 sky130_fd_sc_hd__o31a_1 _14945_ (.A1(net544),
    .A2(net207),
    .A3(_04758_),
    .B1(_05959_),
    .X(_05960_));
 sky130_fd_sc_hd__mux4_1 _14946_ (.A0(net643),
    .A1(net634),
    .A2(net626),
    .A3(net618),
    .S0(net616),
    .S1(net598),
    .X(_05961_));
 sky130_fd_sc_hd__nand2_1 _14947_ (.A(net152),
    .B(_05961_),
    .Y(_05962_));
 sky130_fd_sc_hd__nor3_1 _14948_ (.A(net287),
    .B(_07987_),
    .C(_02819_),
    .Y(_05963_));
 sky130_fd_sc_hd__nor2_1 _14949_ (.A(_00287_),
    .B(_02817_),
    .Y(_05964_));
 sky130_fd_sc_hd__a211o_1 _14950_ (.A1(net289),
    .A2(_05964_),
    .B1(_05963_),
    .C1(net150),
    .X(_05966_));
 sky130_fd_sc_hd__mux2_1 _14951_ (.A0(_05962_),
    .A1(_05966_),
    .S(net296),
    .X(_05967_));
 sky130_fd_sc_hd__nor2_1 _14952_ (.A(_00574_),
    .B(_02815_),
    .Y(_05968_));
 sky130_fd_sc_hd__a21o_1 _14953_ (.A1(net284),
    .A2(net713),
    .B1(_00974_),
    .X(_05969_));
 sky130_fd_sc_hd__nor2_1 _14954_ (.A(net594),
    .B(_05969_),
    .Y(_05970_));
 sky130_fd_sc_hd__a211o_1 _14955_ (.A1(net597),
    .A2(_05968_),
    .B1(_05970_),
    .C1(net150),
    .X(_05971_));
 sky130_fd_sc_hd__nor2_1 _14956_ (.A(_01225_),
    .B(_02848_),
    .Y(_05972_));
 sky130_fd_sc_hd__a21o_1 _14957_ (.A1(net284),
    .A2(net750),
    .B1(_01451_),
    .X(_05973_));
 sky130_fd_sc_hd__nor2_1 _14958_ (.A(net601),
    .B(_05973_),
    .Y(_05974_));
 sky130_fd_sc_hd__a211o_1 _14959_ (.A1(net601),
    .A2(_05972_),
    .B1(_05974_),
    .C1(net150),
    .X(_05975_));
 sky130_fd_sc_hd__mux2_1 _14960_ (.A0(_05971_),
    .A1(_05975_),
    .S(net298),
    .X(_05977_));
 sky130_fd_sc_hd__mux2_4 _14961_ (.A0(_05967_),
    .A1(_05977_),
    .S(net302),
    .X(_05978_));
 sky130_fd_sc_hd__nor2_1 _14962_ (.A(net309),
    .B(net241),
    .Y(_05979_));
 sky130_fd_sc_hd__or2_4 _14963_ (.A(net309),
    .B(net241),
    .X(_05980_));
 sky130_fd_sc_hd__o211ai_4 _14964_ (.A1(_05978_),
    .A2(_05980_),
    .B1(_05940_),
    .C1(_05960_),
    .Y(_05981_));
 sky130_fd_sc_hd__o22a_1 _14965_ (.A1(_03302_),
    .A2(_05880_),
    .B1(_05922_),
    .B2(_05981_),
    .X(_08684_));
 sky130_fd_sc_hd__a21o_1 _14966_ (.A1(net311),
    .A2(_05902_),
    .B1(_05885_),
    .X(_05982_));
 sky130_fd_sc_hd__or4_1 _14967_ (.A(net818),
    .B(net828),
    .C(_05903_),
    .D(_05913_),
    .X(_05983_));
 sky130_fd_sc_hd__a21o_4 _14968_ (.A1(_05982_),
    .A2(_05983_),
    .B1(net314),
    .X(_05984_));
 sky130_fd_sc_hd__a21oi_2 _14969_ (.A1(_05909_),
    .A2(_05984_),
    .B1(net282),
    .Y(_05985_));
 sky130_fd_sc_hd__a21o_4 _14970_ (.A1(_05909_),
    .A2(_05984_),
    .B1(net282),
    .X(_05987_));
 sky130_fd_sc_hd__a21o_1 _14971_ (.A1(\sel_op[1] ),
    .A2(_02584_),
    .B1(_05885_),
    .X(_05988_));
 sky130_fd_sc_hd__a21o_1 _14972_ (.A1(_05883_),
    .A2(_05988_),
    .B1(net312),
    .X(_05989_));
 sky130_fd_sc_hd__a21oi_4 _14973_ (.A1(_05895_),
    .A2(_05989_),
    .B1(net292),
    .Y(_05990_));
 sky130_fd_sc_hd__inv_2 _14974_ (.A(net145),
    .Y(_05991_));
 sky130_fd_sc_hd__or4_4 _14975_ (.A(_05901_),
    .B(_05920_),
    .C(_05987_),
    .D(_05991_),
    .X(_05992_));
 sky130_fd_sc_hd__a22o_1 _14976_ (.A1(net154),
    .A2(net148),
    .B1(net145),
    .B2(net153),
    .X(_05993_));
 sky130_fd_sc_hd__and3_2 _14977_ (.A(net280),
    .B(_05992_),
    .C(_05993_),
    .X(_05994_));
 sky130_fd_sc_hd__nor2_1 _14978_ (.A(_07313_),
    .B(_02610_),
    .Y(_05995_));
 sky130_fd_sc_hd__nor2_1 _14979_ (.A(net289),
    .B(_02606_),
    .Y(_05996_));
 sky130_fd_sc_hd__a211o_1 _14980_ (.A1(net289),
    .A2(_05995_),
    .B1(_05996_),
    .C1(net150),
    .X(_05998_));
 sky130_fd_sc_hd__nor2_1 _14981_ (.A(_07302_),
    .B(_02608_),
    .Y(_05999_));
 sky130_fd_sc_hd__nor3_1 _14982_ (.A(net594),
    .B(_00144_),
    .C(_02603_),
    .Y(_06000_));
 sky130_fd_sc_hd__a211o_1 _14983_ (.A1(net597),
    .A2(_05999_),
    .B1(_06000_),
    .C1(net150),
    .X(_06001_));
 sky130_fd_sc_hd__mux2_1 _14984_ (.A0(_05998_),
    .A1(_06001_),
    .S(net296),
    .X(_06002_));
 sky130_fd_sc_hd__mux4_1 _14985_ (.A0(net710),
    .A1(net697),
    .A2(net688),
    .A3(net679),
    .S0(net609),
    .S1(net596),
    .X(_06003_));
 sky130_fd_sc_hd__nand2_1 _14986_ (.A(net152),
    .B(_06003_),
    .Y(_06004_));
 sky130_fd_sc_hd__mux4_1 _14987_ (.A0(net745),
    .A1(net736),
    .A2(net724),
    .A3(net719),
    .S0(net607),
    .S1(net596),
    .X(_06005_));
 sky130_fd_sc_hd__nand2_1 _14988_ (.A(net152),
    .B(_06005_),
    .Y(_06006_));
 sky130_fd_sc_hd__mux2_1 _14989_ (.A0(_06004_),
    .A1(_06006_),
    .S(net297),
    .X(_06007_));
 sky130_fd_sc_hd__mux2_2 _14990_ (.A0(_06002_),
    .A1(_06007_),
    .S(net301),
    .X(_06009_));
 sky130_fd_sc_hd__mux4_1 _14991_ (.A0(net862),
    .A1(net852),
    .A2(net845),
    .A3(net838),
    .S0(net607),
    .S1(net596),
    .X(_06010_));
 sky130_fd_sc_hd__nand2_1 _14992_ (.A(net152),
    .B(_06010_),
    .Y(_06011_));
 sky130_fd_sc_hd__mux4_1 _14993_ (.A0(net902),
    .A1(net900),
    .A2(net886),
    .A3(net875),
    .S0(net609),
    .S1(net597),
    .X(_06012_));
 sky130_fd_sc_hd__nand2_1 _14994_ (.A(net152),
    .B(_06012_),
    .Y(_06013_));
 sky130_fd_sc_hd__mux2_1 _14995_ (.A0(_06011_),
    .A1(_06013_),
    .S(net297),
    .X(_06014_));
 sky130_fd_sc_hd__mux4_1 _14996_ (.A0(net829),
    .A1(net819),
    .A2(net807),
    .A3(net793),
    .S0(net607),
    .S1(net597),
    .X(_06015_));
 sky130_fd_sc_hd__mux4_1 _14997_ (.A0(net783),
    .A1(net771),
    .A2(net760),
    .A3(net750),
    .S0(net607),
    .S1(net596),
    .X(_06016_));
 sky130_fd_sc_hd__nand2_1 _14998_ (.A(net152),
    .B(_06015_),
    .Y(_06017_));
 sky130_fd_sc_hd__nand2_1 _14999_ (.A(net152),
    .B(_06016_),
    .Y(_06018_));
 sky130_fd_sc_hd__mux2_1 _15000_ (.A0(_06017_),
    .A1(_06018_),
    .S(net584),
    .X(_06020_));
 sky130_fd_sc_hd__mux2_1 _15001_ (.A0(_06014_),
    .A1(_06020_),
    .S(net576),
    .X(_06021_));
 sky130_fd_sc_hd__a21o_1 _15002_ (.A1(net605),
    .A2(net272),
    .B1(net282),
    .X(_06022_));
 sky130_fd_sc_hd__or3_2 _15003_ (.A(net292),
    .B(net906),
    .C(net269),
    .X(_06023_));
 sky130_fd_sc_hd__a21oi_1 _15004_ (.A1(_06022_),
    .A2(_06023_),
    .B1(_05956_),
    .Y(_06024_));
 sky130_fd_sc_hd__a311o_1 _15005_ (.A1(_05956_),
    .A2(_06022_),
    .A3(_06023_),
    .B1(_06024_),
    .C1(net228),
    .X(_06025_));
 sky130_fd_sc_hd__o21ai_1 _15006_ (.A1(_02448_),
    .A2(_05794_),
    .B1(_02446_),
    .Y(_06026_));
 sky130_fd_sc_hd__o311a_1 _15007_ (.A1(_02446_),
    .A2(_02448_),
    .A3(_05794_),
    .B1(net254),
    .C1(_06026_),
    .X(_06027_));
 sky130_fd_sc_hd__or2_1 _15008_ (.A(net905),
    .B(net914),
    .X(_06028_));
 sky130_fd_sc_hd__a32o_1 _15009_ (.A1(_05849_),
    .A2(_05851_),
    .A3(_06028_),
    .B1(net234),
    .B2(net905),
    .X(_06029_));
 sky130_fd_sc_hd__a22o_1 _15010_ (.A1(net615),
    .A2(net905),
    .B1(net915),
    .B2(net603),
    .X(_06031_));
 sky130_fd_sc_hd__and3_1 _15011_ (.A(_02470_),
    .B(net261),
    .C(_06031_),
    .X(_06032_));
 sky130_fd_sc_hd__a2111o_1 _15012_ (.A1(_05795_),
    .A2(net240),
    .B1(_06029_),
    .C1(_06032_),
    .D1(net242),
    .X(_06033_));
 sky130_fd_sc_hd__a211oi_2 _15013_ (.A1(_02448_),
    .A2(net237),
    .B1(_06027_),
    .C1(_06033_),
    .Y(_06034_));
 sky130_fd_sc_hd__o21ai_1 _15014_ (.A1(_05980_),
    .A2(_06009_),
    .B1(_06025_),
    .Y(_06035_));
 sky130_fd_sc_hd__o31a_1 _15015_ (.A1(net559),
    .A2(net210),
    .A3(_02649_),
    .B1(_06034_),
    .X(_06036_));
 sky130_fd_sc_hd__o21ai_1 _15016_ (.A1(net202),
    .A2(_06021_),
    .B1(_06036_),
    .Y(_06037_));
 sky130_fd_sc_hd__o32a_1 _15017_ (.A1(_05994_),
    .A2(_06035_),
    .A3(_06037_),
    .B1(_05880_),
    .B2(net282),
    .X(_08695_));
 sky130_fd_sc_hd__o32a_2 _15018_ (.A1(net818),
    .A2(_05903_),
    .A3(_05913_),
    .B1(_05911_),
    .B2(_05885_),
    .X(_06038_));
 sky130_fd_sc_hd__o22ai_4 _15019_ (.A1(net858),
    .A2(_05907_),
    .B1(_06038_),
    .B2(net313),
    .Y(_06039_));
 sky130_fd_sc_hd__and2_1 _15020_ (.A(net899),
    .B(_06039_),
    .X(_06041_));
 sky130_fd_sc_hd__nand2_4 _15021_ (.A(net899),
    .B(_06039_),
    .Y(_06042_));
 sky130_fd_sc_hd__a22o_2 _15022_ (.A1(net148),
    .A2(net145),
    .B1(net144),
    .B2(net154),
    .X(_06043_));
 sky130_fd_sc_hd__or4_4 _15023_ (.A(_05901_),
    .B(_05987_),
    .C(_05991_),
    .D(_06042_),
    .X(_06044_));
 sky130_fd_sc_hd__a21oi_4 _15024_ (.A1(_05882_),
    .A2(_05886_),
    .B1(net312),
    .Y(_06045_));
 sky130_fd_sc_hd__nor2_2 _15025_ (.A(net533),
    .B(_05897_),
    .Y(_06046_));
 sky130_fd_sc_hd__o21a_4 _15026_ (.A1(_06045_),
    .A2(_06046_),
    .B1(net591),
    .X(_06047_));
 sky130_fd_sc_hd__o21ai_4 _15027_ (.A1(_06045_),
    .A2(_06046_),
    .B1(net591),
    .Y(_06048_));
 sky130_fd_sc_hd__or2_4 _15028_ (.A(_05992_),
    .B(_06048_),
    .X(_06049_));
 sky130_fd_sc_hd__o21ai_4 _15029_ (.A1(_05920_),
    .A2(_06048_),
    .B1(_05992_),
    .Y(_06050_));
 sky130_fd_sc_hd__nand4_4 _15030_ (.A(_06043_),
    .B(_06044_),
    .C(_06049_),
    .D(_06050_),
    .Y(_06052_));
 sky130_fd_sc_hd__a22o_1 _15031_ (.A1(_06043_),
    .A2(_06044_),
    .B1(_06049_),
    .B2(_06050_),
    .X(_06053_));
 sky130_fd_sc_hd__o211ai_4 _15032_ (.A1(_05899_),
    .A2(_02826_),
    .B1(net152),
    .C1(net289),
    .Y(_06054_));
 sky130_fd_sc_hd__mux4_1 _15033_ (.A0(net661),
    .A1(net653),
    .A2(net643),
    .A3(net634),
    .S0(net609),
    .S1(net596),
    .X(_06055_));
 sky130_fd_sc_hd__nand2_1 _15034_ (.A(net152),
    .B(_06055_),
    .Y(_06056_));
 sky130_fd_sc_hd__mux2_1 _15035_ (.A0(_06054_),
    .A1(_06056_),
    .S(net297),
    .X(_06057_));
 sky130_fd_sc_hd__mux2_1 _15036_ (.A0(_05964_),
    .A1(_05968_),
    .S(net289),
    .X(_06058_));
 sky130_fd_sc_hd__or2_2 _15037_ (.A(_05924_),
    .B(_06058_),
    .X(_06059_));
 sky130_fd_sc_hd__nor2_1 _15038_ (.A(net289),
    .B(_05969_),
    .Y(_06060_));
 sky130_fd_sc_hd__a211o_1 _15039_ (.A1(net289),
    .A2(_05972_),
    .B1(_06060_),
    .C1(net150),
    .X(_06061_));
 sky130_fd_sc_hd__mux4_2 _15040_ (.A0(_06054_),
    .A1(_06056_),
    .A2(_06059_),
    .A3(_06061_),
    .S0(net297),
    .S1(net302),
    .X(_06063_));
 sky130_fd_sc_hd__a21o_1 _15041_ (.A1(net592),
    .A2(net276),
    .B1(_03280_),
    .X(_06064_));
 sky130_fd_sc_hd__or3_4 _15042_ (.A(net299),
    .B(net899),
    .C(net269),
    .X(_06065_));
 sky130_fd_sc_hd__a21bo_2 _15043_ (.A1(_05956_),
    .A2(_06023_),
    .B1_N(_06022_),
    .X(_06066_));
 sky130_fd_sc_hd__a21oi_2 _15044_ (.A1(_06064_),
    .A2(_06065_),
    .B1(_06066_),
    .Y(_06067_));
 sky130_fd_sc_hd__a31o_1 _15045_ (.A1(_06064_),
    .A2(_06065_),
    .A3(_06066_),
    .B1(net228),
    .X(_06068_));
 sky130_fd_sc_hd__a21oi_1 _15046_ (.A1(net906),
    .A2(net914),
    .B1(net898),
    .Y(_06069_));
 sky130_fd_sc_hd__a22o_1 _15047_ (.A1(_02386_),
    .A2(net237),
    .B1(net231),
    .B2(net898),
    .X(_06070_));
 sky130_fd_sc_hd__a211oi_1 _15048_ (.A1(_05793_),
    .A2(net240),
    .B1(_06070_),
    .C1(net242),
    .Y(_06071_));
 sky130_fd_sc_hd__o31a_1 _15049_ (.A1(_05850_),
    .A2(_05852_),
    .A3(_06069_),
    .B1(_06071_),
    .X(_06072_));
 sky130_fd_sc_hd__a22o_1 _15050_ (.A1(_02387_),
    .A2(_05793_),
    .B1(_05795_),
    .B2(_05796_),
    .X(_06074_));
 sky130_fd_sc_hd__or3b_1 _15051_ (.A(_05797_),
    .B(net253),
    .C_N(_06074_),
    .X(_06075_));
 sky130_fd_sc_hd__a21oi_1 _15052_ (.A1(_02446_),
    .A2(_02448_),
    .B1(_02449_),
    .Y(_06076_));
 sky130_fd_sc_hd__a31o_1 _15053_ (.A1(_02445_),
    .A2(_02446_),
    .A3(_02448_),
    .B1(_06076_),
    .X(_06077_));
 sky130_fd_sc_hd__o211a_1 _15054_ (.A1(net256),
    .A2(_06077_),
    .B1(_06075_),
    .C1(_06072_),
    .X(_06078_));
 sky130_fd_sc_hd__o31a_1 _15055_ (.A1(net558),
    .A2(net210),
    .A3(_02857_),
    .B1(_06078_),
    .X(_06079_));
 sky130_fd_sc_hd__nor2_1 _15056_ (.A(net289),
    .B(_05973_),
    .Y(_06080_));
 sky130_fd_sc_hd__a211o_1 _15057_ (.A1(net289),
    .A2(_05925_),
    .B1(_06080_),
    .C1(net150),
    .X(_06081_));
 sky130_fd_sc_hd__mux4_1 _15058_ (.A0(net819),
    .A1(net806),
    .A2(net793),
    .A3(net783),
    .S0(net610),
    .S1(net600),
    .X(_06082_));
 sky130_fd_sc_hd__nand2_1 _15059_ (.A(net151),
    .B(_06082_),
    .Y(_06083_));
 sky130_fd_sc_hd__mux4_1 _15060_ (.A0(net855),
    .A1(net845),
    .A2(net838),
    .A3(net829),
    .S0(net610),
    .S1(net600),
    .X(_06085_));
 sky130_fd_sc_hd__nand2_1 _15061_ (.A(net151),
    .B(_06085_),
    .Y(_06086_));
 sky130_fd_sc_hd__mux4_1 _15062_ (.A0(net898),
    .A1(net886),
    .A2(net875),
    .A3(net868),
    .S0(net610),
    .S1(net600),
    .X(_06087_));
 sky130_fd_sc_hd__nand2_1 _15063_ (.A(net151),
    .B(_06087_),
    .Y(_06088_));
 sky130_fd_sc_hd__mux4_2 _15064_ (.A0(_06081_),
    .A1(_06083_),
    .A2(_06086_),
    .A3(_06088_),
    .S0(net299),
    .S1(net303),
    .X(_06089_));
 sky130_fd_sc_hd__o22ai_4 _15065_ (.A1(_05980_),
    .A2(_06063_),
    .B1(_06067_),
    .B2(_06068_),
    .Y(_06090_));
 sky130_fd_sc_hd__o21ai_4 _15066_ (.A1(net202),
    .A2(_06089_),
    .B1(_06079_),
    .Y(_06091_));
 sky130_fd_sc_hd__a31o_1 _15067_ (.A1(net280),
    .A2(_06052_),
    .A3(_06053_),
    .B1(_06091_),
    .X(_06092_));
 sky130_fd_sc_hd__o22a_1 _15068_ (.A1(_03280_),
    .A2(_05880_),
    .B1(_06090_),
    .B2(_06092_),
    .X(_08706_));
 sky130_fd_sc_hd__and2_1 _15069_ (.A(net451),
    .B(net311),
    .X(_06093_));
 sky130_fd_sc_hd__o22a_1 _15070_ (.A1(_02587_),
    .A2(_05881_),
    .B1(_05885_),
    .B2(_06093_),
    .X(_06095_));
 sky130_fd_sc_hd__nor2_2 _15071_ (.A(net312),
    .B(_06095_),
    .Y(_06096_));
 sky130_fd_sc_hd__o21a_2 _15072_ (.A1(_05896_),
    .A2(_06096_),
    .B1(net579),
    .X(_06097_));
 sky130_fd_sc_hd__o21ai_4 _15073_ (.A1(_05896_),
    .A2(_06096_),
    .B1(net579),
    .Y(_06098_));
 sky130_fd_sc_hd__nand2_8 _15074_ (.A(net153),
    .B(net140),
    .Y(_06099_));
 sky130_fd_sc_hd__and2_1 _15075_ (.A(net763),
    .B(\sel_op[1] ),
    .X(_06100_));
 sky130_fd_sc_hd__o22a_1 _15076_ (.A1(_05903_),
    .A2(_05913_),
    .B1(_06100_),
    .B2(_05885_),
    .X(_06101_));
 sky130_fd_sc_hd__nor2_4 _15077_ (.A(net313),
    .B(_06101_),
    .Y(_06102_));
 sky130_fd_sc_hd__o21a_4 _15078_ (.A1(_05908_),
    .A2(_06102_),
    .B1(net889),
    .X(_06103_));
 sky130_fd_sc_hd__o21ai_4 _15079_ (.A1(_05908_),
    .A2(_06102_),
    .B1(net889),
    .Y(_06104_));
 sky130_fd_sc_hd__nand2_4 _15080_ (.A(net145),
    .B(_06103_),
    .Y(_06106_));
 sky130_fd_sc_hd__nor2_2 _15081_ (.A(_05901_),
    .B(net138),
    .Y(_06107_));
 sky130_fd_sc_hd__and3_1 _15082_ (.A(net145),
    .B(net144),
    .C(_06107_),
    .X(_06108_));
 sky130_fd_sc_hd__a22o_1 _15083_ (.A1(net145),
    .A2(net143),
    .B1(_06103_),
    .B2(net154),
    .X(_06109_));
 sky130_fd_sc_hd__o31a_1 _15084_ (.A1(_05901_),
    .A2(_06042_),
    .A3(_06106_),
    .B1(_06109_),
    .X(_06110_));
 sky130_fd_sc_hd__nand2b_1 _15085_ (.A_N(_06099_),
    .B(_06110_),
    .Y(_06111_));
 sky130_fd_sc_hd__a21o_1 _15086_ (.A1(net153),
    .A2(_06097_),
    .B1(_06110_),
    .X(_06112_));
 sky130_fd_sc_hd__nand2_1 _15087_ (.A(_06111_),
    .B(_06112_),
    .Y(_06113_));
 sky130_fd_sc_hd__nand2_1 _15088_ (.A(net148),
    .B(net141),
    .Y(_06114_));
 sky130_fd_sc_hd__mux2_1 _15089_ (.A0(net141),
    .A1(_06114_),
    .S(_06044_),
    .X(_06115_));
 sky130_fd_sc_hd__nand2_1 _15090_ (.A(_06113_),
    .B(_06115_),
    .Y(_06117_));
 sky130_fd_sc_hd__or2_4 _15091_ (.A(_06113_),
    .B(_06115_),
    .X(_06118_));
 sky130_fd_sc_hd__nand2_2 _15092_ (.A(_06117_),
    .B(_06118_),
    .Y(_06119_));
 sky130_fd_sc_hd__nand2_2 _15093_ (.A(_06049_),
    .B(_06052_),
    .Y(_06120_));
 sky130_fd_sc_hd__xor2_4 _15094_ (.A(_06119_),
    .B(_06120_),
    .X(_06121_));
 sky130_fd_sc_hd__or3b_4 _15095_ (.A(net150),
    .B(net596),
    .C_N(_02606_),
    .X(_06122_));
 sky130_fd_sc_hd__mux2_1 _15096_ (.A0(_05995_),
    .A1(_05999_),
    .S(net289),
    .X(_06123_));
 sky130_fd_sc_hd__or2_2 _15097_ (.A(net150),
    .B(_06123_),
    .X(_06124_));
 sky130_fd_sc_hd__mux2_1 _15098_ (.A0(_06122_),
    .A1(_06124_),
    .S(net299),
    .X(_06125_));
 sky130_fd_sc_hd__mux4_1 _15099_ (.A0(net688),
    .A1(net678),
    .A2(net669),
    .A3(net661),
    .S0(net609),
    .S1(net596),
    .X(_06126_));
 sky130_fd_sc_hd__nand2_1 _15100_ (.A(net152),
    .B(_06126_),
    .Y(_06128_));
 sky130_fd_sc_hd__mux4_1 _15101_ (.A0(net724),
    .A1(net719),
    .A2(net705),
    .A3(net701),
    .S0(net610),
    .S1(net601),
    .X(_06129_));
 sky130_fd_sc_hd__nand2_1 _15102_ (.A(_05923_),
    .B(_06129_),
    .Y(_06130_));
 sky130_fd_sc_hd__mux2_1 _15103_ (.A0(_06128_),
    .A1(_06130_),
    .S(net299),
    .X(_06131_));
 sky130_fd_sc_hd__mux2_1 _15104_ (.A0(_06125_),
    .A1(_06131_),
    .S(net303),
    .X(_06132_));
 sky130_fd_sc_hd__o21a_1 _15105_ (.A1(_02471_),
    .A2(_02473_),
    .B1(net261),
    .X(_06133_));
 sky130_fd_sc_hd__nand2_1 _15106_ (.A(_02474_),
    .B(_06133_),
    .Y(_06134_));
 sky130_fd_sc_hd__a21o_1 _15107_ (.A1(_02265_),
    .A2(_05792_),
    .B1(_05798_),
    .X(_06135_));
 sky130_fd_sc_hd__nand2_1 _15108_ (.A(net254),
    .B(_06135_),
    .Y(_06136_));
 sky130_fd_sc_hd__a31o_1 _15109_ (.A1(_02265_),
    .A2(_05792_),
    .A3(_05798_),
    .B1(_06136_),
    .X(_06137_));
 sky130_fd_sc_hd__nor2_1 _15110_ (.A(net886),
    .B(_05852_),
    .Y(_06139_));
 sky130_fd_sc_hd__a22o_1 _15111_ (.A1(_02264_),
    .A2(net237),
    .B1(net231),
    .B2(net886),
    .X(_06140_));
 sky130_fd_sc_hd__a211oi_1 _15112_ (.A1(_05792_),
    .A2(net240),
    .B1(_06140_),
    .C1(net242),
    .Y(_06141_));
 sky130_fd_sc_hd__o311a_1 _15113_ (.A1(net249),
    .A2(_05853_),
    .A3(_06139_),
    .B1(_06141_),
    .C1(_06137_),
    .X(_06142_));
 sky130_fd_sc_hd__o31a_1 _15114_ (.A1(net558),
    .A2(net210),
    .A3(_03022_),
    .B1(_06142_),
    .X(_06143_));
 sky130_fd_sc_hd__o21ai_2 _15115_ (.A1(net303),
    .A2(net270),
    .B1(net890),
    .Y(_06144_));
 sky130_fd_sc_hd__or3_1 _15116_ (.A(net303),
    .B(net890),
    .C(net270),
    .X(_06145_));
 sky130_fd_sc_hd__nand2_1 _15117_ (.A(_06144_),
    .B(_06145_),
    .Y(_06146_));
 sky130_fd_sc_hd__a21boi_4 _15118_ (.A1(_06065_),
    .A2(_06066_),
    .B1_N(_06064_),
    .Y(_06147_));
 sky130_fd_sc_hd__nor2_1 _15119_ (.A(_06146_),
    .B(_06147_),
    .Y(_06148_));
 sky130_fd_sc_hd__a21o_1 _15120_ (.A1(_06146_),
    .A2(_06147_),
    .B1(net228),
    .X(_06150_));
 sky130_fd_sc_hd__a211o_1 _15121_ (.A1(net286),
    .A2(net760),
    .B1(_01547_),
    .C1(net601),
    .X(_06151_));
 sky130_fd_sc_hd__o311a_1 _15122_ (.A1(net292),
    .A2(_01337_),
    .A3(_02636_),
    .B1(net151),
    .C1(_06151_),
    .X(_06152_));
 sky130_fd_sc_hd__inv_2 _15123_ (.A(_06152_),
    .Y(_06153_));
 sky130_fd_sc_hd__mux4_1 _15124_ (.A0(net806),
    .A1(net793),
    .A2(net783),
    .A3(net771),
    .S0(net615),
    .S1(net601),
    .X(_06154_));
 sky130_fd_sc_hd__nand2_1 _15125_ (.A(net151),
    .B(_06154_),
    .Y(_06155_));
 sky130_fd_sc_hd__nand2_1 _15126_ (.A(net587),
    .B(_06152_),
    .Y(_06156_));
 sky130_fd_sc_hd__o21ai_1 _15127_ (.A1(net587),
    .A2(_06155_),
    .B1(_06156_),
    .Y(_06157_));
 sky130_fd_sc_hd__mux4_1 _15128_ (.A0(net845),
    .A1(net838),
    .A2(net829),
    .A3(net816),
    .S0(net615),
    .S1(net605),
    .X(_06158_));
 sky130_fd_sc_hd__mux4_1 _15129_ (.A0(net886),
    .A1(net875),
    .A2(net868),
    .A3(net855),
    .S0(net615),
    .S1(net601),
    .X(_06159_));
 sky130_fd_sc_hd__mux2_1 _15130_ (.A0(_06158_),
    .A1(_06159_),
    .S(net299),
    .X(_06161_));
 sky130_fd_sc_hd__nand2_1 _15131_ (.A(net151),
    .B(_06158_),
    .Y(_06162_));
 sky130_fd_sc_hd__o21a_1 _15132_ (.A1(_06148_),
    .A2(_06150_),
    .B1(_06134_),
    .X(_06163_));
 sky130_fd_sc_hd__o211a_1 _15133_ (.A1(net277),
    .A2(_06121_),
    .B1(_06143_),
    .C1(_06163_),
    .X(_06164_));
 sky130_fd_sc_hd__a31o_1 _15134_ (.A1(net303),
    .A2(net151),
    .A3(_06161_),
    .B1(net558),
    .X(_06165_));
 sky130_fd_sc_hd__a21oi_1 _15135_ (.A1(net577),
    .A2(_06157_),
    .B1(_06165_),
    .Y(_06166_));
 sky130_fd_sc_hd__a211o_1 _15136_ (.A1(net559),
    .A2(_06132_),
    .B1(_06166_),
    .C1(net241),
    .X(_06167_));
 sky130_fd_sc_hd__a22oi_1 _15137_ (.A1(net890),
    .A2(net242),
    .B1(_06164_),
    .B2(_06167_),
    .Y(_08709_));
 sky130_fd_sc_hd__nor2_2 _15138_ (.A(_05987_),
    .B(_06098_),
    .Y(_06168_));
 sky130_fd_sc_hd__nor3_2 _15139_ (.A(net310),
    .B(\sel_op[3] ),
    .C(net311),
    .Y(_06169_));
 sky130_fd_sc_hd__nor2_2 _15140_ (.A(net314),
    .B(_06169_),
    .Y(_06171_));
 sky130_fd_sc_hd__or2_4 _15141_ (.A(net314),
    .B(_06169_),
    .X(_06172_));
 sky130_fd_sc_hd__o21a_1 _15142_ (.A1(net451),
    .A2(net461),
    .B1(net310),
    .X(_06173_));
 sky130_fd_sc_hd__or3_4 _15143_ (.A(net313),
    .B(net268),
    .C(_06173_),
    .X(_06174_));
 sky130_fd_sc_hd__a2111o_1 _15144_ (.A1(_02585_),
    .A2(_05885_),
    .B1(net268),
    .C1(_06173_),
    .D1(net312),
    .X(_06175_));
 sky130_fd_sc_hd__a21o_4 _15145_ (.A1(_05894_),
    .A2(_06175_),
    .B1(net309),
    .X(_06176_));
 sky130_fd_sc_hd__or3_4 _15146_ (.A(_03302_),
    .B(_05918_),
    .C(net200),
    .X(_06177_));
 sky130_fd_sc_hd__nor4_4 _15147_ (.A(net310),
    .B(\sel_op[3] ),
    .C(net311),
    .D(net314),
    .Y(_06178_));
 sky130_fd_sc_hd__nand2_8 _15148_ (.A(_03335_),
    .B(net268),
    .Y(_06179_));
 sky130_fd_sc_hd__o41a_1 _15149_ (.A1(net763),
    .A2(net774),
    .A3(net785),
    .A4(net796),
    .B1(\sel_op[2] ),
    .X(_06180_));
 sky130_fd_sc_hd__o32a_1 _15150_ (.A1(_05902_),
    .A2(_05904_),
    .A3(_05905_),
    .B1(_06180_),
    .B2(net313),
    .X(_06182_));
 sky130_fd_sc_hd__and3b_4 _15151_ (.A_N(_06182_),
    .B(net878),
    .C(net227),
    .X(_06183_));
 sky130_fd_sc_hd__or3b_4 _15152_ (.A(net266),
    .B(_06182_),
    .C_N(net878),
    .X(_06184_));
 sky130_fd_sc_hd__a211o_4 _15153_ (.A1(_05890_),
    .A2(_05898_),
    .B1(_06184_),
    .C1(net286),
    .X(_06185_));
 sky130_fd_sc_hd__or2_2 _15154_ (.A(_06177_),
    .B(_06185_),
    .X(_06186_));
 sky130_fd_sc_hd__xor2_4 _15155_ (.A(_06177_),
    .B(_06185_),
    .X(_06187_));
 sky130_fd_sc_hd__nand2b_2 _15156_ (.A_N(_06106_),
    .B(_06187_),
    .Y(_06188_));
 sky130_fd_sc_hd__xnor2_4 _15157_ (.A(_06106_),
    .B(_06187_),
    .Y(_06189_));
 sky130_fd_sc_hd__nand2_2 _15158_ (.A(_06168_),
    .B(_06189_),
    .Y(_06190_));
 sky130_fd_sc_hd__xnor2_1 _15159_ (.A(_06168_),
    .B(_06189_),
    .Y(_06191_));
 sky130_fd_sc_hd__or2_2 _15160_ (.A(_06111_),
    .B(_06191_),
    .X(_06193_));
 sky130_fd_sc_hd__nand2_1 _15161_ (.A(_06111_),
    .B(_06191_),
    .Y(_06194_));
 sky130_fd_sc_hd__nand2_4 _15162_ (.A(_06193_),
    .B(_06194_),
    .Y(_06195_));
 sky130_fd_sc_hd__a21o_1 _15163_ (.A1(net144),
    .A2(net141),
    .B1(_06108_),
    .X(_06196_));
 sky130_fd_sc_hd__nand2_2 _15164_ (.A(net141),
    .B(_06108_),
    .Y(_06197_));
 sky130_fd_sc_hd__nand2_4 _15165_ (.A(_06196_),
    .B(_06197_),
    .Y(_06198_));
 sky130_fd_sc_hd__xnor2_4 _15166_ (.A(_06195_),
    .B(_06198_),
    .Y(_06199_));
 sky130_fd_sc_hd__o21ai_4 _15167_ (.A1(_06044_),
    .A2(_06048_),
    .B1(_06118_),
    .Y(_06200_));
 sky130_fd_sc_hd__nand2b_1 _15168_ (.A_N(_06199_),
    .B(_06200_),
    .Y(_06201_));
 sky130_fd_sc_hd__xnor2_4 _15169_ (.A(_06199_),
    .B(_06200_),
    .Y(_06202_));
 sky130_fd_sc_hd__and3_2 _15170_ (.A(_06117_),
    .B(_06118_),
    .C(_06120_),
    .X(_06204_));
 sky130_fd_sc_hd__xnor2_2 _15171_ (.A(_06202_),
    .B(_06204_),
    .Y(_06205_));
 sky130_fd_sc_hd__a21oi_1 _15172_ (.A1(_02474_),
    .A2(_02477_),
    .B1(net257),
    .Y(_06206_));
 sky130_fd_sc_hd__nand2_1 _15173_ (.A(_02478_),
    .B(_06206_),
    .Y(_06207_));
 sky130_fd_sc_hd__o21ai_1 _15174_ (.A1(net309),
    .A2(net269),
    .B1(net878),
    .Y(_06208_));
 sky130_fd_sc_hd__or3_2 _15175_ (.A(net309),
    .B(net875),
    .C(net269),
    .X(_06209_));
 sky130_fd_sc_hd__o21ai_2 _15176_ (.A1(_06146_),
    .A2(_06147_),
    .B1(_06144_),
    .Y(_06210_));
 sky130_fd_sc_hd__a21oi_1 _15177_ (.A1(_06208_),
    .A2(_06209_),
    .B1(_06210_),
    .Y(_06211_));
 sky130_fd_sc_hd__a311o_1 _15178_ (.A1(_06208_),
    .A2(_06209_),
    .A3(_06210_),
    .B1(_06211_),
    .C1(net228),
    .X(_06212_));
 sky130_fd_sc_hd__mux2_1 _15179_ (.A0(_05966_),
    .A1(_05971_),
    .S(net298),
    .X(_06213_));
 sky130_fd_sc_hd__or2_2 _15180_ (.A(net584),
    .B(_05962_),
    .X(_06215_));
 sky130_fd_sc_hd__o22a_1 _15181_ (.A1(_03689_),
    .A2(_05962_),
    .B1(_06213_),
    .B2(net575),
    .X(_06216_));
 sky130_fd_sc_hd__o21ai_1 _15182_ (.A1(_02116_),
    .A2(_05791_),
    .B1(_05799_),
    .Y(_06217_));
 sky130_fd_sc_hd__o311a_1 _15183_ (.A1(_02116_),
    .A2(_05791_),
    .A3(_05799_),
    .B1(net254),
    .C1(_06217_),
    .X(_06218_));
 sky130_fd_sc_hd__a2bb2o_1 _15184_ (.A1_N(_05791_),
    .A2_N(_05942_),
    .B1(net231),
    .B2(net876),
    .X(_06219_));
 sky130_fd_sc_hd__a21oi_1 _15185_ (.A1(net875),
    .A2(_05853_),
    .B1(net249),
    .Y(_06220_));
 sky130_fd_sc_hd__o21a_1 _15186_ (.A1(net875),
    .A2(_05853_),
    .B1(_06220_),
    .X(_06221_));
 sky130_fd_sc_hd__a2111o_1 _15187_ (.A1(_02116_),
    .A2(net237),
    .B1(_06219_),
    .C1(_06221_),
    .D1(net242),
    .X(_06222_));
 sky130_fd_sc_hd__nor2_1 _15188_ (.A(_06218_),
    .B(_06222_),
    .Y(_06223_));
 sky130_fd_sc_hd__a21oi_1 _15189_ (.A1(net151),
    .A2(_05934_),
    .B1(net592),
    .Y(_06224_));
 sky130_fd_sc_hd__a211o_1 _15190_ (.A1(net592),
    .A2(_05930_),
    .B1(_06224_),
    .C1(net576),
    .X(_06226_));
 sky130_fd_sc_hd__mux2_1 _15191_ (.A0(_05928_),
    .A1(_05975_),
    .S(net592),
    .X(_06227_));
 sky130_fd_sc_hd__o21a_1 _15192_ (.A1(net304),
    .A2(_06227_),
    .B1(_06226_),
    .X(_06228_));
 sky130_fd_sc_hd__o221a_1 _15193_ (.A1(_05980_),
    .A2(_06216_),
    .B1(_06228_),
    .B2(net202),
    .C1(_06223_),
    .X(_06229_));
 sky130_fd_sc_hd__o311a_1 _15194_ (.A1(net544),
    .A2(net207),
    .A3(_03194_),
    .B1(_06212_),
    .C1(_06229_),
    .X(_06230_));
 sky130_fd_sc_hd__o211a_2 _15195_ (.A1(net277),
    .A2(_06205_),
    .B1(_06207_),
    .C1(_06230_),
    .X(_06231_));
 sky130_fd_sc_hd__a21oi_1 _15196_ (.A1(net879),
    .A2(net244),
    .B1(_06231_),
    .Y(_08710_));
 sky130_fd_sc_hd__nand2_4 _15197_ (.A(net144),
    .B(net140),
    .Y(_06232_));
 sky130_fd_sc_hd__a21o_2 _15198_ (.A1(\sel_op[2] ),
    .A2(_02584_),
    .B1(_06172_),
    .X(_06233_));
 sky130_fd_sc_hd__a21boi_4 _15199_ (.A1(_05893_),
    .A2(_06233_),
    .B1_N(net547),
    .Y(_06234_));
 sky130_fd_sc_hd__a21bo_4 _15200_ (.A1(_05893_),
    .A2(_06233_),
    .B1_N(net547),
    .X(_06236_));
 sky130_fd_sc_hd__nand2_4 _15201_ (.A(net153),
    .B(net136),
    .Y(_06237_));
 sky130_fd_sc_hd__a211o_4 _15202_ (.A1(_05909_),
    .A2(_05984_),
    .B1(net200),
    .C1(net282),
    .X(_06238_));
 sky130_fd_sc_hd__a21o_2 _15203_ (.A1(_05885_),
    .A2(_05913_),
    .B1(net313),
    .X(_06239_));
 sky130_fd_sc_hd__or3b_4 _15204_ (.A(net764),
    .B(net774),
    .C_N(net312),
    .X(_06240_));
 sky130_fd_sc_hd__nor2_2 _15205_ (.A(_05912_),
    .B(_06240_),
    .Y(_06241_));
 sky130_fd_sc_hd__and2_1 _15206_ (.A(_03269_),
    .B(_06241_),
    .X(_06242_));
 sky130_fd_sc_hd__or3_4 _15207_ (.A(_03335_),
    .B(_05902_),
    .C(_05904_),
    .X(_06243_));
 sky130_fd_sc_hd__or4_4 _15208_ (.A(net828),
    .B(_03335_),
    .C(_05902_),
    .D(_05904_),
    .X(_06244_));
 sky130_fd_sc_hd__a21boi_4 _15209_ (.A1(_06239_),
    .A2(_06244_),
    .B1_N(net867),
    .Y(_06245_));
 sky130_fd_sc_hd__a21bo_4 _15210_ (.A1(_06239_),
    .A2(_06244_),
    .B1_N(net867),
    .X(_06247_));
 sky130_fd_sc_hd__a211oi_4 _15211_ (.A1(_05890_),
    .A2(_05898_),
    .B1(net196),
    .C1(net286),
    .Y(_06248_));
 sky130_fd_sc_hd__nor2_1 _15212_ (.A(net200),
    .B(net196),
    .Y(_06249_));
 sky130_fd_sc_hd__and3_1 _15213_ (.A(net154),
    .B(net148),
    .C(_06249_),
    .X(_06250_));
 sky130_fd_sc_hd__xnor2_4 _15214_ (.A(_06238_),
    .B(_06248_),
    .Y(_06251_));
 sky130_fd_sc_hd__nand2_2 _15215_ (.A(net145),
    .B(net198),
    .Y(_06252_));
 sky130_fd_sc_hd__xor2_4 _15216_ (.A(_06251_),
    .B(_06252_),
    .X(_06253_));
 sky130_fd_sc_hd__or2_4 _15217_ (.A(_06237_),
    .B(_06253_),
    .X(_06254_));
 sky130_fd_sc_hd__xor2_4 _15218_ (.A(_06237_),
    .B(_06253_),
    .X(_06255_));
 sky130_fd_sc_hd__nand2b_4 _15219_ (.A_N(_06232_),
    .B(_06255_),
    .Y(_06256_));
 sky130_fd_sc_hd__xnor2_4 _15220_ (.A(_06232_),
    .B(_06255_),
    .Y(_06258_));
 sky130_fd_sc_hd__xnor2_4 _15221_ (.A(_06190_),
    .B(_06258_),
    .Y(_06259_));
 sky130_fd_sc_hd__nand2_2 _15222_ (.A(_06186_),
    .B(_06188_),
    .Y(_06260_));
 sky130_fd_sc_hd__nand2_4 _15223_ (.A(net141),
    .B(_06103_),
    .Y(_06261_));
 sky130_fd_sc_hd__a21o_4 _15224_ (.A1(_06186_),
    .A2(_06188_),
    .B1(_06261_),
    .X(_06262_));
 sky130_fd_sc_hd__xnor2_4 _15225_ (.A(_06260_),
    .B(_06261_),
    .Y(_06263_));
 sky130_fd_sc_hd__xnor2_2 _15226_ (.A(_06259_),
    .B(_06263_),
    .Y(_06264_));
 sky130_fd_sc_hd__o21a_1 _15227_ (.A1(_06195_),
    .A2(_06198_),
    .B1(_06193_),
    .X(_06265_));
 sky130_fd_sc_hd__xnor2_1 _15228_ (.A(_06264_),
    .B(_06265_),
    .Y(_06266_));
 sky130_fd_sc_hd__or2_1 _15229_ (.A(_06197_),
    .B(_06266_),
    .X(_06267_));
 sky130_fd_sc_hd__nand2_1 _15230_ (.A(_06197_),
    .B(_06266_),
    .Y(_06269_));
 sky130_fd_sc_hd__nand2_1 _15231_ (.A(_06267_),
    .B(_06269_),
    .Y(_06270_));
 sky130_fd_sc_hd__a21boi_2 _15232_ (.A1(_06202_),
    .A2(_06204_),
    .B1_N(_06201_),
    .Y(_06271_));
 sky130_fd_sc_hd__or2_4 _15233_ (.A(_06270_),
    .B(_06271_),
    .X(_06272_));
 sky130_fd_sc_hd__a21oi_2 _15234_ (.A1(_06270_),
    .A2(_06271_),
    .B1(net279),
    .Y(_06273_));
 sky130_fd_sc_hd__nand3_1 _15235_ (.A(_02469_),
    .B(_02476_),
    .C(_02478_),
    .Y(_06274_));
 sky130_fd_sc_hd__a21o_1 _15236_ (.A1(_02476_),
    .A2(_02478_),
    .B1(_02469_),
    .X(_06275_));
 sky130_fd_sc_hd__a21bo_1 _15237_ (.A1(net544),
    .A2(net272),
    .B1_N(net868),
    .X(_06276_));
 sky130_fd_sc_hd__or3b_2 _15238_ (.A(net868),
    .B(net269),
    .C_N(net544),
    .X(_06277_));
 sky130_fd_sc_hd__a21bo_2 _15239_ (.A1(_06209_),
    .A2(_06210_),
    .B1_N(_06208_),
    .X(_06278_));
 sky130_fd_sc_hd__a21o_1 _15240_ (.A1(_06276_),
    .A2(_06277_),
    .B1(_06278_),
    .X(_06280_));
 sky130_fd_sc_hd__nand3_1 _15241_ (.A(_06276_),
    .B(_06277_),
    .C(_06278_),
    .Y(_06281_));
 sky130_fd_sc_hd__and3_1 _15242_ (.A(net230),
    .B(_06280_),
    .C(_06281_),
    .X(_06282_));
 sky130_fd_sc_hd__o21ai_1 _15243_ (.A1(_02060_),
    .A2(_05789_),
    .B1(_05800_),
    .Y(_06283_));
 sky130_fd_sc_hd__or3_1 _15244_ (.A(_02060_),
    .B(_05789_),
    .C(_05800_),
    .X(_06284_));
 sky130_fd_sc_hd__mux2_1 _15245_ (.A0(_06001_),
    .A1(_06004_),
    .S(net297),
    .X(_06285_));
 sky130_fd_sc_hd__o22a_1 _15246_ (.A1(_03689_),
    .A2(_05998_),
    .B1(_06285_),
    .B2(net566),
    .X(_06286_));
 sky130_fd_sc_hd__a31o_1 _15247_ (.A1(net875),
    .A2(net886),
    .A3(_05852_),
    .B1(net868),
    .X(_06287_));
 sky130_fd_sc_hd__and3b_1 _15248_ (.A_N(_05854_),
    .B(_06287_),
    .C(_05849_),
    .X(_06288_));
 sky130_fd_sc_hd__a2bb2o_1 _15249_ (.A1_N(_05789_),
    .A2_N(_05942_),
    .B1(net231),
    .B2(net865),
    .X(_06289_));
 sky130_fd_sc_hd__a211o_1 _15250_ (.A1(_02060_),
    .A2(net237),
    .B1(_06289_),
    .C1(net242),
    .X(_06291_));
 sky130_fd_sc_hd__a31o_1 _15251_ (.A1(net254),
    .A2(_06283_),
    .A3(_06284_),
    .B1(_06291_),
    .X(_06292_));
 sky130_fd_sc_hd__or2_2 _15252_ (.A(net585),
    .B(_05998_),
    .X(_06293_));
 sky130_fd_sc_hd__mux2_1 _15253_ (.A0(_06006_),
    .A1(_06018_),
    .S(net297),
    .X(_06294_));
 sky130_fd_sc_hd__mux2_1 _15254_ (.A0(_06011_),
    .A1(_06017_),
    .S(net584),
    .X(_06295_));
 sky130_fd_sc_hd__mux4_1 _15255_ (.A0(_06285_),
    .A1(_06293_),
    .A2(_06295_),
    .A3(_06294_),
    .S0(net566),
    .S1(net308),
    .X(_06296_));
 sky130_fd_sc_hd__o32a_1 _15256_ (.A1(net558),
    .A2(net209),
    .A3(_03360_),
    .B1(net241),
    .B2(_06296_),
    .X(_06297_));
 sky130_fd_sc_hd__or4b_4 _15257_ (.A(_06282_),
    .B(_06288_),
    .C(_06292_),
    .D_N(_06297_),
    .X(_06298_));
 sky130_fd_sc_hd__a31o_2 _15258_ (.A1(net261),
    .A2(_06274_),
    .A3(_06275_),
    .B1(_06298_),
    .X(_06299_));
 sky130_fd_sc_hd__a21oi_4 _15259_ (.A1(_06272_),
    .A2(_06273_),
    .B1(_06299_),
    .Y(_06300_));
 sky130_fd_sc_hd__a21oi_4 _15260_ (.A1(net867),
    .A2(net247),
    .B1(_06300_),
    .Y(_08711_));
 sky130_fd_sc_hd__nand2_4 _15261_ (.A(net140),
    .B(_06103_),
    .Y(_06302_));
 sky130_fd_sc_hd__or4_4 _15262_ (.A(net490),
    .B(net500),
    .C(_03335_),
    .D(_02586_),
    .X(_06303_));
 sky130_fd_sc_hd__a21boi_4 _15263_ (.A1(_06174_),
    .A2(_06303_),
    .B1_N(net532),
    .Y(_06304_));
 sky130_fd_sc_hd__a21bo_4 _15264_ (.A1(_06174_),
    .A2(_06303_),
    .B1_N(net533),
    .X(_06305_));
 sky130_fd_sc_hd__a211o_4 _15265_ (.A1(_05909_),
    .A2(_05984_),
    .B1(_06305_),
    .C1(net282),
    .X(_06306_));
 sky130_fd_sc_hd__or3_4 _15266_ (.A(_05920_),
    .B(_06236_),
    .C(_06306_),
    .X(_06307_));
 sky130_fd_sc_hd__a22o_1 _15267_ (.A1(net148),
    .A2(net136),
    .B1(net194),
    .B2(net153),
    .X(_06308_));
 sky130_fd_sc_hd__nand2_4 _15268_ (.A(_06307_),
    .B(_06308_),
    .Y(_06309_));
 sky130_fd_sc_hd__o21a_1 _15269_ (.A1(net763),
    .A2(net774),
    .B1(\sel_op[2] ),
    .X(_06310_));
 sky130_fd_sc_hd__or3_4 _15270_ (.A(net313),
    .B(net268),
    .C(_06310_),
    .X(_06312_));
 sky130_fd_sc_hd__a21boi_4 _15271_ (.A1(_06243_),
    .A2(_06312_),
    .B1_N(net858),
    .Y(_06313_));
 sky130_fd_sc_hd__a21bo_1 _15272_ (.A1(_06243_),
    .A2(_06312_),
    .B1_N(net858),
    .X(_06314_));
 sky130_fd_sc_hd__nor2_1 _15273_ (.A(net200),
    .B(net192),
    .Y(_06315_));
 sky130_fd_sc_hd__or3b_4 _15274_ (.A(_03280_),
    .B(net200),
    .C_N(_06039_),
    .X(_06316_));
 sky130_fd_sc_hd__a211o_4 _15275_ (.A1(_05890_),
    .A2(_05898_),
    .B1(net192),
    .C1(net286),
    .X(_06317_));
 sky130_fd_sc_hd__nor2_1 _15276_ (.A(_06316_),
    .B(_06317_),
    .Y(_06318_));
 sky130_fd_sc_hd__xor2_4 _15277_ (.A(_06316_),
    .B(_06317_),
    .X(_06319_));
 sky130_fd_sc_hd__nand2_2 _15278_ (.A(net145),
    .B(_06245_),
    .Y(_06320_));
 sky130_fd_sc_hd__xor2_4 _15279_ (.A(_06319_),
    .B(_06320_),
    .X(_06321_));
 sky130_fd_sc_hd__nor2_4 _15280_ (.A(_06309_),
    .B(_06321_),
    .Y(_06323_));
 sky130_fd_sc_hd__xnor2_4 _15281_ (.A(_06309_),
    .B(_06321_),
    .Y(_06324_));
 sky130_fd_sc_hd__nor2_1 _15282_ (.A(_06254_),
    .B(_06324_),
    .Y(_06325_));
 sky130_fd_sc_hd__xnor2_4 _15283_ (.A(_06254_),
    .B(_06324_),
    .Y(_06326_));
 sky130_fd_sc_hd__or2_4 _15284_ (.A(_06302_),
    .B(_06326_),
    .X(_06327_));
 sky130_fd_sc_hd__xnor2_4 _15285_ (.A(_06302_),
    .B(_06326_),
    .Y(_06328_));
 sky130_fd_sc_hd__nor2_1 _15286_ (.A(_06256_),
    .B(_06328_),
    .Y(_06329_));
 sky130_fd_sc_hd__xor2_4 _15287_ (.A(_06256_),
    .B(_06328_),
    .X(_06330_));
 sky130_fd_sc_hd__a31o_4 _15288_ (.A1(net145),
    .A2(net198),
    .A3(_06251_),
    .B1(_06250_),
    .X(_06331_));
 sky130_fd_sc_hd__nand2_2 _15289_ (.A(net141),
    .B(net198),
    .Y(_06332_));
 sky130_fd_sc_hd__and3_1 _15290_ (.A(net141),
    .B(net198),
    .C(_06331_),
    .X(_06334_));
 sky130_fd_sc_hd__xnor2_4 _15291_ (.A(_06331_),
    .B(_06332_),
    .Y(_06335_));
 sky130_fd_sc_hd__xnor2_4 _15292_ (.A(_06330_),
    .B(_06335_),
    .Y(_06336_));
 sky130_fd_sc_hd__a32o_4 _15293_ (.A1(_06168_),
    .A2(_06189_),
    .A3(_06258_),
    .B1(_06259_),
    .B2(_06263_),
    .X(_06337_));
 sky130_fd_sc_hd__nand2b_1 _15294_ (.A_N(_06336_),
    .B(_06337_),
    .Y(_06338_));
 sky130_fd_sc_hd__xor2_4 _15295_ (.A(_06336_),
    .B(_06337_),
    .X(_06339_));
 sky130_fd_sc_hd__xnor2_4 _15296_ (.A(_06262_),
    .B(_06339_),
    .Y(_06340_));
 sky130_fd_sc_hd__o21a_2 _15297_ (.A1(_06264_),
    .A2(_06265_),
    .B1(_06267_),
    .X(_06341_));
 sky130_fd_sc_hd__nor2_1 _15298_ (.A(_06340_),
    .B(_06341_),
    .Y(_06342_));
 sky130_fd_sc_hd__xnor2_4 _15299_ (.A(_06340_),
    .B(_06341_),
    .Y(_06343_));
 sky130_fd_sc_hd__a21oi_1 _15300_ (.A1(_06272_),
    .A2(_06343_),
    .B1(net279),
    .Y(_06345_));
 sky130_fd_sc_hd__o21ai_2 _15301_ (.A1(_06272_),
    .A2(_06343_),
    .B1(_06345_),
    .Y(_06346_));
 sky130_fd_sc_hd__or2_1 _15302_ (.A(_02479_),
    .B(_02483_),
    .X(_06347_));
 sky130_fd_sc_hd__nand2_1 _15303_ (.A(_02484_),
    .B(_06347_),
    .Y(_06348_));
 sky130_fd_sc_hd__a21boi_1 _15304_ (.A1(net534),
    .A2(net272),
    .B1_N(net855),
    .Y(_06349_));
 sky130_fd_sc_hd__and3b_1 _15305_ (.A_N(net855),
    .B(net272),
    .C(net534),
    .X(_06350_));
 sky130_fd_sc_hd__a21boi_2 _15306_ (.A1(_06277_),
    .A2(_06278_),
    .B1_N(_06276_),
    .Y(_06351_));
 sky130_fd_sc_hd__or3_1 _15307_ (.A(_06349_),
    .B(_06350_),
    .C(_06351_),
    .X(_06352_));
 sky130_fd_sc_hd__o21a_1 _15308_ (.A1(_06349_),
    .A2(_06350_),
    .B1(_06351_),
    .X(_06353_));
 sky130_fd_sc_hd__or3b_1 _15309_ (.A(_06353_),
    .B(net228),
    .C_N(_06352_),
    .X(_06354_));
 sky130_fd_sc_hd__o21a_1 _15310_ (.A1(_01662_),
    .A2(_05788_),
    .B1(_05802_),
    .X(_06356_));
 sky130_fd_sc_hd__or3b_1 _15311_ (.A(net253),
    .B(_06356_),
    .C_N(_05803_),
    .X(_06357_));
 sky130_fd_sc_hd__mux2_2 _15312_ (.A0(_06056_),
    .A1(_06059_),
    .S(net297),
    .X(_06358_));
 sky130_fd_sc_hd__o22ai_4 _15313_ (.A1(_03689_),
    .A2(_06054_),
    .B1(_06358_),
    .B2(net575),
    .Y(_06359_));
 sky130_fd_sc_hd__nor2_1 _15314_ (.A(net855),
    .B(_05854_),
    .Y(_06360_));
 sky130_fd_sc_hd__or3_1 _15315_ (.A(net249),
    .B(_05855_),
    .C(_06360_),
    .X(_06361_));
 sky130_fd_sc_hd__o2bb2a_1 _15316_ (.A1_N(net857),
    .A2_N(net231),
    .B1(_05942_),
    .B2(_05788_),
    .X(_06362_));
 sky130_fd_sc_hd__o211a_1 _15317_ (.A1(_01663_),
    .A2(net235),
    .B1(_06362_),
    .C1(_05880_),
    .X(_06363_));
 sky130_fd_sc_hd__o311a_1 _15318_ (.A1(net558),
    .A2(net210),
    .A3(_03527_),
    .B1(_06361_),
    .C1(_06363_),
    .X(_06364_));
 sky130_fd_sc_hd__mux4_1 _15319_ (.A0(_06061_),
    .A1(_06081_),
    .A2(_06083_),
    .A3(_06086_),
    .S0(net299),
    .S1(net303),
    .X(_06365_));
 sky130_fd_sc_hd__o2bb2a_1 _15320_ (.A1_N(_05979_),
    .A2_N(_06359_),
    .B1(_06365_),
    .B2(net202),
    .X(_06367_));
 sky130_fd_sc_hd__and4_2 _15321_ (.A(_06354_),
    .B(_06357_),
    .C(_06364_),
    .D(_06367_),
    .X(_06368_));
 sky130_fd_sc_hd__o211a_2 _15322_ (.A1(net256),
    .A2(_06348_),
    .B1(_06368_),
    .C1(_06346_),
    .X(_06369_));
 sky130_fd_sc_hd__a21oi_1 _15323_ (.A1(net859),
    .A2(net244),
    .B1(_06369_),
    .Y(_08712_));
 sky130_fd_sc_hd__nand2_4 _15324_ (.A(net140),
    .B(net198),
    .Y(_06370_));
 sky130_fd_sc_hd__a211o_2 _15325_ (.A1(net452),
    .A2(net310),
    .B1(net312),
    .C1(net268),
    .X(_06371_));
 sky130_fd_sc_hd__a21oi_4 _15326_ (.A1(_05891_),
    .A2(_06371_),
    .B1(_03182_),
    .Y(_06372_));
 sky130_fd_sc_hd__a21o_1 _15327_ (.A1(_05891_),
    .A2(_06371_),
    .B1(_03182_),
    .X(_06373_));
 sky130_fd_sc_hd__a211o_1 _15328_ (.A1(_05909_),
    .A2(_05984_),
    .B1(net190),
    .C1(_03291_),
    .X(_06374_));
 sky130_fd_sc_hd__or3_4 _15329_ (.A(_03302_),
    .B(_05918_),
    .C(net190),
    .X(_06375_));
 sky130_fd_sc_hd__nor2_1 _15330_ (.A(_06306_),
    .B(_06375_),
    .Y(_06377_));
 sky130_fd_sc_hd__xor2_4 _15331_ (.A(_06306_),
    .B(_06375_),
    .X(_06378_));
 sky130_fd_sc_hd__nand2_2 _15332_ (.A(net144),
    .B(net136),
    .Y(_06379_));
 sky130_fd_sc_hd__and3_1 _15333_ (.A(net144),
    .B(net136),
    .C(_06378_),
    .X(_06380_));
 sky130_fd_sc_hd__xor2_4 _15334_ (.A(_06378_),
    .B(_06379_),
    .X(_06381_));
 sky130_fd_sc_hd__nor2_1 _15335_ (.A(_06307_),
    .B(_06381_),
    .Y(_06382_));
 sky130_fd_sc_hd__nand2_1 _15336_ (.A(_06307_),
    .B(_06381_),
    .Y(_06383_));
 sky130_fd_sc_hd__xnor2_4 _15337_ (.A(_06307_),
    .B(_06381_),
    .Y(_06384_));
 sky130_fd_sc_hd__a21oi_2 _15338_ (.A1(net763),
    .A2(net310),
    .B1(_06172_),
    .Y(_06385_));
 sky130_fd_sc_hd__o21ai_4 _15339_ (.A1(_06242_),
    .A2(_06385_),
    .B1(net848),
    .Y(_06386_));
 sky130_fd_sc_hd__o22a_4 _15340_ (.A1(net138),
    .A2(net200),
    .B1(net135),
    .B2(_05901_),
    .X(_06388_));
 sky130_fd_sc_hd__nor2_8 _15341_ (.A(net200),
    .B(net135),
    .Y(_06389_));
 sky130_fd_sc_hd__nand2_1 _15342_ (.A(_06107_),
    .B(_06389_),
    .Y(_06390_));
 sky130_fd_sc_hd__a21oi_4 _15343_ (.A1(_06107_),
    .A2(_06389_),
    .B1(_06388_),
    .Y(_06391_));
 sky130_fd_sc_hd__nand2_4 _15344_ (.A(net146),
    .B(net193),
    .Y(_06392_));
 sky130_fd_sc_hd__xnor2_4 _15345_ (.A(_06391_),
    .B(_06392_),
    .Y(_06393_));
 sky130_fd_sc_hd__xnor2_4 _15346_ (.A(_06384_),
    .B(_06393_),
    .Y(_06394_));
 sky130_fd_sc_hd__nand2_2 _15347_ (.A(_06323_),
    .B(_06394_),
    .Y(_06395_));
 sky130_fd_sc_hd__xnor2_4 _15348_ (.A(_06323_),
    .B(_06394_),
    .Y(_06396_));
 sky130_fd_sc_hd__nor2_4 _15349_ (.A(_06370_),
    .B(_06396_),
    .Y(_06397_));
 sky130_fd_sc_hd__xnor2_4 _15350_ (.A(_06370_),
    .B(_06396_),
    .Y(_06399_));
 sky130_fd_sc_hd__or2_2 _15351_ (.A(_06327_),
    .B(_06399_),
    .X(_06400_));
 sky130_fd_sc_hd__xnor2_4 _15352_ (.A(_06327_),
    .B(_06399_),
    .Y(_06401_));
 sky130_fd_sc_hd__a31o_1 _15353_ (.A1(net145),
    .A2(_06245_),
    .A3(_06319_),
    .B1(_06318_),
    .X(_06402_));
 sky130_fd_sc_hd__nand2_2 _15354_ (.A(_06325_),
    .B(_06402_),
    .Y(_06403_));
 sky130_fd_sc_hd__or2_2 _15355_ (.A(_06325_),
    .B(_06402_),
    .X(_06404_));
 sky130_fd_sc_hd__nand2_4 _15356_ (.A(_06403_),
    .B(_06404_),
    .Y(_06405_));
 sky130_fd_sc_hd__nand2_4 _15357_ (.A(net141),
    .B(_06245_),
    .Y(_06406_));
 sky130_fd_sc_hd__xnor2_4 _15358_ (.A(_06405_),
    .B(_06406_),
    .Y(_06407_));
 sky130_fd_sc_hd__xor2_4 _15359_ (.A(_06401_),
    .B(_06407_),
    .X(_06408_));
 sky130_fd_sc_hd__a21oi_2 _15360_ (.A1(_06330_),
    .A2(_06335_),
    .B1(_06329_),
    .Y(_06410_));
 sky130_fd_sc_hd__nand2b_1 _15361_ (.A_N(_06410_),
    .B(_06408_),
    .Y(_06411_));
 sky130_fd_sc_hd__xnor2_2 _15362_ (.A(_06408_),
    .B(_06410_),
    .Y(_06412_));
 sky130_fd_sc_hd__xnor2_1 _15363_ (.A(_06334_),
    .B(_06412_),
    .Y(_06413_));
 sky130_fd_sc_hd__o21ai_2 _15364_ (.A1(_06262_),
    .A2(_06339_),
    .B1(_06338_),
    .Y(_06414_));
 sky130_fd_sc_hd__and2b_1 _15365_ (.A_N(_06413_),
    .B(_06414_),
    .X(_06415_));
 sky130_fd_sc_hd__nand2b_1 _15366_ (.A_N(_06414_),
    .B(_06413_),
    .Y(_06416_));
 sky130_fd_sc_hd__nand2b_1 _15367_ (.A_N(_06415_),
    .B(_06416_),
    .Y(_06417_));
 sky130_fd_sc_hd__o21bai_4 _15368_ (.A1(_06272_),
    .A2(_06343_),
    .B1_N(_06342_),
    .Y(_06418_));
 sky130_fd_sc_hd__xnor2_2 _15369_ (.A(_06417_),
    .B(_06418_),
    .Y(_06419_));
 sky130_fd_sc_hd__a21o_1 _15370_ (.A1(_02482_),
    .A2(_02485_),
    .B1(_02488_),
    .X(_06421_));
 sky130_fd_sc_hd__a211o_1 _15371_ (.A1(_02484_),
    .A2(_06421_),
    .B1(net257),
    .C1(_02486_),
    .X(_06422_));
 sky130_fd_sc_hd__o21a_1 _15372_ (.A1(_03182_),
    .A2(net269),
    .B1(net845),
    .X(_06423_));
 sky130_fd_sc_hd__and3b_1 _15373_ (.A_N(net849),
    .B(net272),
    .C(net523),
    .X(_06424_));
 sky130_fd_sc_hd__or2_1 _15374_ (.A(_06423_),
    .B(_06424_),
    .X(_06425_));
 sky130_fd_sc_hd__o21ba_1 _15375_ (.A1(_06350_),
    .A2(_06351_),
    .B1_N(_06349_),
    .X(_06426_));
 sky130_fd_sc_hd__a21oi_1 _15376_ (.A1(_06425_),
    .A2(_06426_),
    .B1(net228),
    .Y(_06427_));
 sky130_fd_sc_hd__o21ai_1 _15377_ (.A1(_06425_),
    .A2(_06426_),
    .B1(_06427_),
    .Y(_06428_));
 sky130_fd_sc_hd__o21a_1 _15378_ (.A1(_01593_),
    .A2(_05787_),
    .B1(_05804_),
    .X(_06429_));
 sky130_fd_sc_hd__a211o_1 _15379_ (.A1(_01594_),
    .A2(_05805_),
    .B1(net253),
    .C1(_06429_),
    .X(_06430_));
 sky130_fd_sc_hd__mux4_1 _15380_ (.A0(_06130_),
    .A1(_06153_),
    .A2(_06155_),
    .A3(_06162_),
    .S0(net299),
    .S1(net303),
    .X(_06432_));
 sky130_fd_sc_hd__nor2_1 _15381_ (.A(net845),
    .B(_05855_),
    .Y(_06433_));
 sky130_fd_sc_hd__o2bb2a_1 _15382_ (.A1_N(net847),
    .A2_N(net231),
    .B1(_05942_),
    .B2(_05787_),
    .X(_06434_));
 sky130_fd_sc_hd__o211a_1 _15383_ (.A1(_01594_),
    .A2(net235),
    .B1(_06434_),
    .C1(_05880_),
    .X(_06435_));
 sky130_fd_sc_hd__mux2_2 _15384_ (.A0(_06124_),
    .A1(_06128_),
    .S(net297),
    .X(_06436_));
 sky130_fd_sc_hd__o22ai_4 _15385_ (.A1(_03689_),
    .A2(_06122_),
    .B1(_06436_),
    .B2(net575),
    .Y(_06437_));
 sky130_fd_sc_hd__nand2_1 _15386_ (.A(_05979_),
    .B(_06437_),
    .Y(_06438_));
 sky130_fd_sc_hd__o311a_1 _15387_ (.A1(net249),
    .A2(_05857_),
    .A3(_06433_),
    .B1(_06435_),
    .C1(_06438_),
    .X(_06439_));
 sky130_fd_sc_hd__o211a_1 _15388_ (.A1(net202),
    .A2(_06432_),
    .B1(_06439_),
    .C1(_06430_),
    .X(_06440_));
 sky130_fd_sc_hd__o311a_1 _15389_ (.A1(net558),
    .A2(net211),
    .A3(_03684_),
    .B1(_06428_),
    .C1(_06440_),
    .X(_06441_));
 sky130_fd_sc_hd__nand2_1 _15390_ (.A(_06422_),
    .B(_06441_),
    .Y(_06443_));
 sky130_fd_sc_hd__a21oi_2 _15391_ (.A1(net280),
    .A2(_06419_),
    .B1(_06443_),
    .Y(_06444_));
 sky130_fd_sc_hd__a21oi_2 _15392_ (.A1(net848),
    .A2(net243),
    .B1(_06444_),
    .Y(_08713_));
 sky130_fd_sc_hd__nand2_2 _15393_ (.A(net478),
    .B(_06172_),
    .Y(_06445_));
 sky130_fd_sc_hd__a21oi_4 _15394_ (.A1(net314),
    .A2(_02584_),
    .B1(net266),
    .Y(_06446_));
 sky130_fd_sc_hd__and3_4 _15395_ (.A(net516),
    .B(_06445_),
    .C(_06446_),
    .X(_06447_));
 sky130_fd_sc_hd__nand3_4 _15396_ (.A(net516),
    .B(_06445_),
    .C(_06446_),
    .Y(_06448_));
 sky130_fd_sc_hd__nand2_8 _15397_ (.A(net197),
    .B(net131),
    .Y(_06449_));
 sky130_fd_sc_hd__nor2_4 _15398_ (.A(_06099_),
    .B(_06449_),
    .Y(_06450_));
 sky130_fd_sc_hd__o22a_1 _15399_ (.A1(_06098_),
    .A2(net196),
    .B1(_06448_),
    .B2(_05920_),
    .X(_06451_));
 sky130_fd_sc_hd__or2_4 _15400_ (.A(_06450_),
    .B(_06451_),
    .X(_06453_));
 sky130_fd_sc_hd__and3_1 _15401_ (.A(net899),
    .B(_06039_),
    .C(net194),
    .X(_06454_));
 sky130_fd_sc_hd__and3_4 _15402_ (.A(net899),
    .B(_06039_),
    .C(_06372_),
    .X(_06455_));
 sky130_fd_sc_hd__and3_1 _15403_ (.A(net148),
    .B(net194),
    .C(_06455_),
    .X(_06456_));
 sky130_fd_sc_hd__xnor2_2 _15404_ (.A(_06374_),
    .B(_06454_),
    .Y(_06457_));
 sky130_fd_sc_hd__nor2_1 _15405_ (.A(net138),
    .B(_06236_),
    .Y(_06458_));
 sky130_fd_sc_hd__xor2_1 _15406_ (.A(_06457_),
    .B(_06458_),
    .X(_06459_));
 sky130_fd_sc_hd__o21a_2 _15407_ (.A1(_06377_),
    .A2(_06380_),
    .B1(_06459_),
    .X(_06460_));
 sky130_fd_sc_hd__or3_4 _15408_ (.A(_06377_),
    .B(_06380_),
    .C(_06459_),
    .X(_06461_));
 sky130_fd_sc_hd__nand2b_4 _15409_ (.A_N(_06460_),
    .B(_06461_),
    .Y(_06462_));
 sky130_fd_sc_hd__o21a_4 _15410_ (.A1(_06171_),
    .A2(_06241_),
    .B1(net837),
    .X(_06464_));
 sky130_fd_sc_hd__o21ai_4 _15411_ (.A1(_06171_),
    .A2(_06241_),
    .B1(net837),
    .Y(_06465_));
 sky130_fd_sc_hd__nor2_4 _15412_ (.A(net200),
    .B(_06184_),
    .Y(_06466_));
 sky130_fd_sc_hd__nand2_4 _15413_ (.A(net154),
    .B(_06464_),
    .Y(_06467_));
 sky130_fd_sc_hd__xor2_4 _15414_ (.A(_06466_),
    .B(_06467_),
    .X(_06468_));
 sky130_fd_sc_hd__or2_4 _15415_ (.A(_05991_),
    .B(net135),
    .X(_06469_));
 sky130_fd_sc_hd__nor2_1 _15416_ (.A(_06468_),
    .B(_06469_),
    .Y(_06470_));
 sky130_fd_sc_hd__xor2_4 _15417_ (.A(_06468_),
    .B(_06469_),
    .X(_06471_));
 sky130_fd_sc_hd__and3b_1 _15418_ (.A_N(_06460_),
    .B(_06461_),
    .C(_06471_),
    .X(_06472_));
 sky130_fd_sc_hd__xor2_4 _15419_ (.A(_06462_),
    .B(_06471_),
    .X(_06473_));
 sky130_fd_sc_hd__a21o_2 _15420_ (.A1(_06383_),
    .A2(_06393_),
    .B1(_06382_),
    .X(_06475_));
 sky130_fd_sc_hd__and2b_2 _15421_ (.A_N(_06473_),
    .B(_06475_),
    .X(_06476_));
 sky130_fd_sc_hd__xor2_4 _15422_ (.A(_06473_),
    .B(_06475_),
    .X(_06477_));
 sky130_fd_sc_hd__nor2_4 _15423_ (.A(_06453_),
    .B(_06477_),
    .Y(_06478_));
 sky130_fd_sc_hd__xor2_4 _15424_ (.A(_06453_),
    .B(_06477_),
    .X(_06479_));
 sky130_fd_sc_hd__nand2_1 _15425_ (.A(_06397_),
    .B(_06479_),
    .Y(_06480_));
 sky130_fd_sc_hd__xor2_4 _15426_ (.A(_06397_),
    .B(_06479_),
    .X(_06481_));
 sky130_fd_sc_hd__o21ai_4 _15427_ (.A1(_06388_),
    .A2(_06392_),
    .B1(_06390_),
    .Y(_06482_));
 sky130_fd_sc_hd__and3_1 _15428_ (.A(_06323_),
    .B(_06394_),
    .C(_06482_),
    .X(_06483_));
 sky130_fd_sc_hd__xnor2_4 _15429_ (.A(_06395_),
    .B(_06482_),
    .Y(_06484_));
 sky130_fd_sc_hd__nand2_2 _15430_ (.A(net142),
    .B(net193),
    .Y(_06486_));
 sky130_fd_sc_hd__xnor2_4 _15431_ (.A(_06484_),
    .B(_06486_),
    .Y(_06487_));
 sky130_fd_sc_hd__nand2_1 _15432_ (.A(_06481_),
    .B(_06487_),
    .Y(_06488_));
 sky130_fd_sc_hd__xor2_4 _15433_ (.A(_06481_),
    .B(_06487_),
    .X(_06489_));
 sky130_fd_sc_hd__o21ai_4 _15434_ (.A1(_06401_),
    .A2(_06407_),
    .B1(_06400_),
    .Y(_06490_));
 sky130_fd_sc_hd__and2_1 _15435_ (.A(_06489_),
    .B(_06490_),
    .X(_06491_));
 sky130_fd_sc_hd__xnor2_4 _15436_ (.A(_06489_),
    .B(_06490_),
    .Y(_06492_));
 sky130_fd_sc_hd__o21ai_4 _15437_ (.A1(_06405_),
    .A2(_06406_),
    .B1(_06403_),
    .Y(_06493_));
 sky130_fd_sc_hd__and2b_1 _15438_ (.A_N(_06492_),
    .B(_06493_),
    .X(_06494_));
 sky130_fd_sc_hd__xor2_4 _15439_ (.A(_06492_),
    .B(_06493_),
    .X(_06495_));
 sky130_fd_sc_hd__a21bo_2 _15440_ (.A1(_06334_),
    .A2(_06412_),
    .B1_N(_06411_),
    .X(_06497_));
 sky130_fd_sc_hd__and2b_1 _15441_ (.A_N(_06495_),
    .B(_06497_),
    .X(_06498_));
 sky130_fd_sc_hd__xnor2_2 _15442_ (.A(_06495_),
    .B(_06497_),
    .Y(_06499_));
 sky130_fd_sc_hd__a21o_2 _15443_ (.A1(_06416_),
    .A2(_06418_),
    .B1(_06415_),
    .X(_06500_));
 sky130_fd_sc_hd__o21ai_1 _15444_ (.A1(_06499_),
    .A2(_06500_),
    .B1(net281),
    .Y(_06501_));
 sky130_fd_sc_hd__a21o_1 _15445_ (.A1(_06499_),
    .A2(_06500_),
    .B1(_06501_),
    .X(_06502_));
 sky130_fd_sc_hd__a211oi_1 _15446_ (.A1(_02467_),
    .A2(_02489_),
    .B1(_02488_),
    .C1(_02486_),
    .Y(_06503_));
 sky130_fd_sc_hd__or2_1 _15447_ (.A(_02490_),
    .B(net257),
    .X(_06504_));
 sky130_fd_sc_hd__a21bo_2 _15448_ (.A1(net516),
    .A2(net272),
    .B1_N(net837),
    .X(_06505_));
 sky130_fd_sc_hd__inv_2 _15449_ (.A(_06505_),
    .Y(_06506_));
 sky130_fd_sc_hd__or3b_2 _15450_ (.A(net837),
    .B(net269),
    .C_N(net516),
    .X(_06508_));
 sky130_fd_sc_hd__o21bai_2 _15451_ (.A1(_06424_),
    .A2(_06426_),
    .B1_N(_06423_),
    .Y(_06509_));
 sky130_fd_sc_hd__a21o_1 _15452_ (.A1(_06505_),
    .A2(_06508_),
    .B1(_06509_),
    .X(_06510_));
 sky130_fd_sc_hd__nand3_1 _15453_ (.A(_06505_),
    .B(_06508_),
    .C(_06509_),
    .Y(_06511_));
 sky130_fd_sc_hd__and3_1 _15454_ (.A(net230),
    .B(_06510_),
    .C(_06511_),
    .X(_06512_));
 sky130_fd_sc_hd__a21o_1 _15455_ (.A1(_01716_),
    .A2(_05786_),
    .B1(_05806_),
    .X(_06513_));
 sky130_fd_sc_hd__or3b_1 _15456_ (.A(_05807_),
    .B(net253),
    .C_N(_06513_),
    .X(_06514_));
 sky130_fd_sc_hd__or3_2 _15457_ (.A(net544),
    .B(_02648_),
    .C(_03690_),
    .X(_06515_));
 sky130_fd_sc_hd__nor2_1 _15458_ (.A(net304),
    .B(_05977_),
    .Y(_06516_));
 sky130_fd_sc_hd__o21ai_1 _15459_ (.A1(net575),
    .A2(_05931_),
    .B1(net309),
    .Y(_06517_));
 sky130_fd_sc_hd__or2_1 _15460_ (.A(net575),
    .B(_05967_),
    .X(_06519_));
 sky130_fd_sc_hd__a21oi_1 _15461_ (.A1(net558),
    .A2(_06519_),
    .B1(net241),
    .Y(_06520_));
 sky130_fd_sc_hd__o21ai_1 _15462_ (.A1(_06516_),
    .A2(_06517_),
    .B1(_06520_),
    .Y(_06521_));
 sky130_fd_sc_hd__nor2_1 _15463_ (.A(net836),
    .B(_05857_),
    .Y(_06522_));
 sky130_fd_sc_hd__a221o_1 _15464_ (.A1(_05786_),
    .A2(net240),
    .B1(net231),
    .B2(net836),
    .C1(net242),
    .X(_06523_));
 sky130_fd_sc_hd__a21oi_1 _15465_ (.A1(_01715_),
    .A2(net237),
    .B1(_06523_),
    .Y(_06524_));
 sky130_fd_sc_hd__o311a_1 _15466_ (.A1(net249),
    .A2(_05858_),
    .A3(_06522_),
    .B1(_06524_),
    .C1(_06521_),
    .X(_06525_));
 sky130_fd_sc_hd__and4b_2 _15467_ (.A_N(_06512_),
    .B(_06514_),
    .C(_06515_),
    .D(_06525_),
    .X(_06526_));
 sky130_fd_sc_hd__o211a_1 _15468_ (.A1(_06503_),
    .A2(_06504_),
    .B1(_06526_),
    .C1(_06502_),
    .X(_06527_));
 sky130_fd_sc_hd__a21oi_2 _15469_ (.A1(net837),
    .A2(net243),
    .B1(_06527_),
    .Y(_08714_));
 sky130_fd_sc_hd__a21o_4 _15470_ (.A1(_06499_),
    .A2(_06500_),
    .B1(_06498_),
    .X(_06529_));
 sky130_fd_sc_hd__and2_4 _15471_ (.A(net507),
    .B(_06446_),
    .X(_06530_));
 sky130_fd_sc_hd__nand2_2 _15472_ (.A(net507),
    .B(_06446_),
    .Y(_06531_));
 sky130_fd_sc_hd__a22o_1 _15473_ (.A1(net148),
    .A2(net131),
    .B1(_06530_),
    .B2(net153),
    .X(_06532_));
 sky130_fd_sc_hd__a211o_4 _15474_ (.A1(_05909_),
    .A2(_05984_),
    .B1(net186),
    .C1(_03291_),
    .X(_06533_));
 sky130_fd_sc_hd__and4_2 _15475_ (.A(net153),
    .B(net148),
    .C(net131),
    .D(_06530_),
    .X(_06534_));
 sky130_fd_sc_hd__inv_2 _15476_ (.A(_06534_),
    .Y(_06535_));
 sky130_fd_sc_hd__or4b_4 _15477_ (.A(_06098_),
    .B(_06534_),
    .C(net192),
    .D_N(_06532_),
    .X(_06536_));
 sky130_fd_sc_hd__a22o_1 _15478_ (.A1(net140),
    .A2(net193),
    .B1(_06532_),
    .B2(_06535_),
    .X(_06537_));
 sky130_fd_sc_hd__nand2_4 _15479_ (.A(_06536_),
    .B(_06537_),
    .Y(_06538_));
 sky130_fd_sc_hd__or3_4 _15480_ (.A(_06099_),
    .B(_06449_),
    .C(_06538_),
    .X(_06540_));
 sky130_fd_sc_hd__xnor2_4 _15481_ (.A(_06450_),
    .B(_06538_),
    .Y(_06541_));
 sky130_fd_sc_hd__o211a_4 _15482_ (.A1(_05908_),
    .A2(_06102_),
    .B1(net194),
    .C1(net889),
    .X(_06542_));
 sky130_fd_sc_hd__nand2_1 _15483_ (.A(_06455_),
    .B(_06542_),
    .Y(_06543_));
 sky130_fd_sc_hd__xnor2_4 _15484_ (.A(_06455_),
    .B(_06542_),
    .Y(_06544_));
 sky130_fd_sc_hd__nand2_4 _15485_ (.A(net198),
    .B(net136),
    .Y(_06545_));
 sky130_fd_sc_hd__xnor2_4 _15486_ (.A(_06544_),
    .B(_06545_),
    .Y(_06546_));
 sky130_fd_sc_hd__a21o_4 _15487_ (.A1(_06457_),
    .A2(_06458_),
    .B1(_06456_),
    .X(_06547_));
 sky130_fd_sc_hd__nand2b_2 _15488_ (.A_N(_06546_),
    .B(_06547_),
    .Y(_06548_));
 sky130_fd_sc_hd__xor2_4 _15489_ (.A(_06546_),
    .B(_06547_),
    .X(_06549_));
 sky130_fd_sc_hd__a21bo_2 _15490_ (.A1(net314),
    .A2(_05902_),
    .B1_N(\ApproximateM_inst.lob_16.lob1.genblk1[9].genblk1.mux.sel ),
    .X(_06551_));
 sky130_fd_sc_hd__nor2_4 _15491_ (.A(net266),
    .B(_06551_),
    .Y(_06552_));
 sky130_fd_sc_hd__or2_4 _15492_ (.A(net266),
    .B(_06551_),
    .X(_06553_));
 sky130_fd_sc_hd__nor2_2 _15493_ (.A(net200),
    .B(_06553_),
    .Y(_06554_));
 sky130_fd_sc_hd__and2_2 _15494_ (.A(_06248_),
    .B(_06554_),
    .X(_06555_));
 sky130_fd_sc_hd__a21oi_2 _15495_ (.A1(net155),
    .A2(net184),
    .B1(_06249_),
    .Y(_06556_));
 sky130_fd_sc_hd__nor2_4 _15496_ (.A(_06555_),
    .B(_06556_),
    .Y(_06557_));
 sky130_fd_sc_hd__nand2_2 _15497_ (.A(net146),
    .B(net188),
    .Y(_06558_));
 sky130_fd_sc_hd__xor2_4 _15498_ (.A(_06557_),
    .B(_06558_),
    .X(_06559_));
 sky130_fd_sc_hd__xor2_2 _15499_ (.A(_06549_),
    .B(_06559_),
    .X(_06560_));
 sky130_fd_sc_hd__o21a_2 _15500_ (.A1(_06460_),
    .A2(_06472_),
    .B1(_06560_),
    .X(_06562_));
 sky130_fd_sc_hd__nor3_2 _15501_ (.A(_06460_),
    .B(_06472_),
    .C(_06560_),
    .Y(_06563_));
 sky130_fd_sc_hd__nor2_4 _15502_ (.A(_06562_),
    .B(_06563_),
    .Y(_06564_));
 sky130_fd_sc_hd__nand2_2 _15503_ (.A(_06541_),
    .B(_06564_),
    .Y(_06565_));
 sky130_fd_sc_hd__xor2_4 _15504_ (.A(_06541_),
    .B(_06564_),
    .X(_06566_));
 sky130_fd_sc_hd__xnor2_2 _15505_ (.A(_06478_),
    .B(_06566_),
    .Y(_06567_));
 sky130_fd_sc_hd__a31o_4 _15506_ (.A1(net155),
    .A2(net188),
    .A3(_06466_),
    .B1(_06470_),
    .X(_06568_));
 sky130_fd_sc_hd__xnor2_4 _15507_ (.A(_06476_),
    .B(_06568_),
    .Y(_06569_));
 sky130_fd_sc_hd__or2_4 _15508_ (.A(_06048_),
    .B(net135),
    .X(_06570_));
 sky130_fd_sc_hd__nor2_1 _15509_ (.A(_06569_),
    .B(_06570_),
    .Y(_06571_));
 sky130_fd_sc_hd__xor2_4 _15510_ (.A(_06569_),
    .B(_06570_),
    .X(_06573_));
 sky130_fd_sc_hd__and2b_1 _15511_ (.A_N(_06567_),
    .B(_06573_),
    .X(_06574_));
 sky130_fd_sc_hd__xor2_2 _15512_ (.A(_06567_),
    .B(_06573_),
    .X(_06575_));
 sky130_fd_sc_hd__a21oi_2 _15513_ (.A1(_06480_),
    .A2(_06488_),
    .B1(_06575_),
    .Y(_06576_));
 sky130_fd_sc_hd__and3_1 _15514_ (.A(_06480_),
    .B(_06488_),
    .C(_06575_),
    .X(_06577_));
 sky130_fd_sc_hd__nor2_1 _15515_ (.A(_06576_),
    .B(_06577_),
    .Y(_06578_));
 sky130_fd_sc_hd__a31oi_4 _15516_ (.A1(net141),
    .A2(net193),
    .A3(_06484_),
    .B1(_06483_),
    .Y(_06579_));
 sky130_fd_sc_hd__and2b_1 _15517_ (.A_N(_06579_),
    .B(_06578_),
    .X(_06580_));
 sky130_fd_sc_hd__xnor2_1 _15518_ (.A(_06578_),
    .B(_06579_),
    .Y(_06581_));
 sky130_fd_sc_hd__o21a_1 _15519_ (.A1(_06491_),
    .A2(_06494_),
    .B1(_06581_),
    .X(_06582_));
 sky130_fd_sc_hd__or3_2 _15520_ (.A(_06491_),
    .B(_06494_),
    .C(_06581_),
    .X(_06584_));
 sky130_fd_sc_hd__nand2b_2 _15521_ (.A_N(_06582_),
    .B(_06584_),
    .Y(_06585_));
 sky130_fd_sc_hd__xor2_4 _15522_ (.A(_06529_),
    .B(_06585_),
    .X(_06586_));
 sky130_fd_sc_hd__or2_1 _15523_ (.A(net277),
    .B(_06586_),
    .X(_06587_));
 sky130_fd_sc_hd__nand3b_1 _15524_ (.A_N(_02419_),
    .B(_02421_),
    .C(_02441_),
    .Y(_06588_));
 sky130_fd_sc_hd__and2_1 _15525_ (.A(_02442_),
    .B(_06588_),
    .X(_06589_));
 sky130_fd_sc_hd__a21o_1 _15526_ (.A1(_02421_),
    .A2(_02465_),
    .B1(_02490_),
    .X(_06590_));
 sky130_fd_sc_hd__a21oi_1 _15527_ (.A1(_06589_),
    .A2(_06590_),
    .B1(net256),
    .Y(_06591_));
 sky130_fd_sc_hd__o21ai_2 _15528_ (.A1(_06589_),
    .A2(_06590_),
    .B1(_06591_),
    .Y(_06592_));
 sky130_fd_sc_hd__a21boi_1 _15529_ (.A1(net507),
    .A2(net272),
    .B1_N(net829),
    .Y(_06593_));
 sky130_fd_sc_hd__or3b_1 _15530_ (.A(net828),
    .B(net269),
    .C_N(net507),
    .X(_06595_));
 sky130_fd_sc_hd__and2b_1 _15531_ (.A_N(_06593_),
    .B(_06595_),
    .X(_06596_));
 sky130_fd_sc_hd__nand2_1 _15532_ (.A(_06505_),
    .B(_06511_),
    .Y(_06597_));
 sky130_fd_sc_hd__xnor2_1 _15533_ (.A(_06596_),
    .B(_06597_),
    .Y(_06598_));
 sky130_fd_sc_hd__a21o_1 _15534_ (.A1(_01414_),
    .A2(_05785_),
    .B1(_05808_),
    .X(_06599_));
 sky130_fd_sc_hd__nand2_1 _15535_ (.A(net254),
    .B(_06599_),
    .Y(_06600_));
 sky130_fd_sc_hd__a31o_1 _15536_ (.A1(_01414_),
    .A2(_05785_),
    .A3(_05808_),
    .B1(_06600_),
    .X(_06601_));
 sky130_fd_sc_hd__or2_2 _15537_ (.A(net575),
    .B(_06002_),
    .X(_06602_));
 sky130_fd_sc_hd__or2_1 _15538_ (.A(net576),
    .B(_06020_),
    .X(_06603_));
 sky130_fd_sc_hd__o211a_1 _15539_ (.A1(net301),
    .A2(_06007_),
    .B1(_06603_),
    .C1(net308),
    .X(_06604_));
 sky130_fd_sc_hd__a211o_1 _15540_ (.A1(net558),
    .A2(_06602_),
    .B1(_06604_),
    .C1(net241),
    .X(_06606_));
 sky130_fd_sc_hd__nor2_1 _15541_ (.A(net827),
    .B(_05858_),
    .Y(_06607_));
 sky130_fd_sc_hd__a221o_1 _15542_ (.A1(_05785_),
    .A2(net240),
    .B1(net231),
    .B2(net827),
    .C1(net242),
    .X(_06608_));
 sky130_fd_sc_hd__o21ba_1 _15543_ (.A1(_01414_),
    .A2(net235),
    .B1_N(_06608_),
    .X(_06609_));
 sky130_fd_sc_hd__o311a_1 _15544_ (.A1(net249),
    .A2(_05859_),
    .A3(_06607_),
    .B1(_06609_),
    .C1(_06606_),
    .X(_06610_));
 sky130_fd_sc_hd__o311a_1 _15545_ (.A1(net544),
    .A2(net207),
    .A3(_03858_),
    .B1(_06601_),
    .C1(_06610_),
    .X(_06611_));
 sky130_fd_sc_hd__o211a_1 _15546_ (.A1(net228),
    .A2(_06598_),
    .B1(_06611_),
    .C1(_06592_),
    .X(_06612_));
 sky130_fd_sc_hd__a22o_1 _15547_ (.A1(net829),
    .A2(net243),
    .B1(_06587_),
    .B2(_06612_),
    .X(_06613_));
 sky130_fd_sc_hd__inv_2 _15548_ (.A(_06613_),
    .Y(_08715_));
 sky130_fd_sc_hd__nor2_4 _15549_ (.A(_06098_),
    .B(net135),
    .Y(_06614_));
 sky130_fd_sc_hd__a21bo_1 _15550_ (.A1(net314),
    .A2(_02583_),
    .B1_N(net500),
    .X(_06616_));
 sky130_fd_sc_hd__nor2_4 _15551_ (.A(net266),
    .B(_06616_),
    .Y(_06617_));
 sky130_fd_sc_hd__or2_1 _15552_ (.A(net267),
    .B(_06616_),
    .X(_06618_));
 sky130_fd_sc_hd__or3_4 _15553_ (.A(_03302_),
    .B(_05918_),
    .C(net181),
    .X(_06619_));
 sky130_fd_sc_hd__nor2_1 _15554_ (.A(_06533_),
    .B(_06619_),
    .Y(_06620_));
 sky130_fd_sc_hd__xor2_4 _15555_ (.A(_06533_),
    .B(_06619_),
    .X(_06621_));
 sky130_fd_sc_hd__nand2_1 _15556_ (.A(net144),
    .B(net131),
    .Y(_06622_));
 sky130_fd_sc_hd__xnor2_2 _15557_ (.A(_06621_),
    .B(_06622_),
    .Y(_06623_));
 sky130_fd_sc_hd__nor2_1 _15558_ (.A(_06534_),
    .B(_06623_),
    .Y(_06624_));
 sky130_fd_sc_hd__nand2_2 _15559_ (.A(_06534_),
    .B(_06623_),
    .Y(_06625_));
 sky130_fd_sc_hd__and2b_4 _15560_ (.A_N(_06624_),
    .B(_06625_),
    .X(_06627_));
 sky130_fd_sc_hd__nand2_1 _15561_ (.A(_06614_),
    .B(_06627_),
    .Y(_06628_));
 sky130_fd_sc_hd__xnor2_4 _15562_ (.A(_06614_),
    .B(_06627_),
    .Y(_06629_));
 sky130_fd_sc_hd__nor2_1 _15563_ (.A(_06536_),
    .B(_06629_),
    .Y(_06630_));
 sky130_fd_sc_hd__xor2_4 _15564_ (.A(_06536_),
    .B(_06629_),
    .X(_06631_));
 sky130_fd_sc_hd__a22o_1 _15565_ (.A1(net198),
    .A2(net194),
    .B1(_06372_),
    .B2(_06103_),
    .X(_06632_));
 sky130_fd_sc_hd__nor2_4 _15566_ (.A(_06184_),
    .B(net190),
    .Y(_06633_));
 sky130_fd_sc_hd__nand2_1 _15567_ (.A(_06542_),
    .B(_06633_),
    .Y(_06634_));
 sky130_fd_sc_hd__and2_2 _15568_ (.A(_06632_),
    .B(_06634_),
    .X(_06635_));
 sky130_fd_sc_hd__nor2_4 _15569_ (.A(_06236_),
    .B(_06247_),
    .Y(_06636_));
 sky130_fd_sc_hd__xor2_4 _15570_ (.A(_06635_),
    .B(_06636_),
    .X(_06638_));
 sky130_fd_sc_hd__o21a_2 _15571_ (.A1(_06544_),
    .A2(_06545_),
    .B1(_06543_),
    .X(_06639_));
 sky130_fd_sc_hd__nand2b_2 _15572_ (.A_N(_06639_),
    .B(_06638_),
    .Y(_06640_));
 sky130_fd_sc_hd__xnor2_4 _15573_ (.A(_06638_),
    .B(_06639_),
    .Y(_06641_));
 sky130_fd_sc_hd__a21oi_4 _15574_ (.A1(net764),
    .A2(net314),
    .B1(net267),
    .Y(_06642_));
 sky130_fd_sc_hd__a21boi_4 _15575_ (.A1(_06172_),
    .A2(_06240_),
    .B1_N(net818),
    .Y(_06643_));
 sky130_fd_sc_hd__a21bo_1 _15576_ (.A1(_06172_),
    .A2(_06240_),
    .B1_N(net818),
    .X(_06644_));
 sky130_fd_sc_hd__nand2_1 _15577_ (.A(net155),
    .B(net178),
    .Y(_06645_));
 sky130_fd_sc_hd__and3_1 _15578_ (.A(net154),
    .B(_06315_),
    .C(net177),
    .X(_06646_));
 sky130_fd_sc_hd__a21oi_2 _15579_ (.A1(net154),
    .A2(net177),
    .B1(_06315_),
    .Y(_06647_));
 sky130_fd_sc_hd__nor2_2 _15580_ (.A(_06646_),
    .B(_06647_),
    .Y(_06649_));
 sky130_fd_sc_hd__nand2_4 _15581_ (.A(net146),
    .B(net184),
    .Y(_06650_));
 sky130_fd_sc_hd__xnor2_4 _15582_ (.A(_06649_),
    .B(_06650_),
    .Y(_06651_));
 sky130_fd_sc_hd__nand2_2 _15583_ (.A(_06641_),
    .B(_06651_),
    .Y(_06652_));
 sky130_fd_sc_hd__xnor2_4 _15584_ (.A(_06641_),
    .B(_06651_),
    .Y(_06653_));
 sky130_fd_sc_hd__o21ai_4 _15585_ (.A1(_06549_),
    .A2(_06559_),
    .B1(_06548_),
    .Y(_06654_));
 sky130_fd_sc_hd__and2b_1 _15586_ (.A_N(_06653_),
    .B(_06654_),
    .X(_06655_));
 sky130_fd_sc_hd__xnor2_4 _15587_ (.A(_06653_),
    .B(_06654_),
    .Y(_06656_));
 sky130_fd_sc_hd__xnor2_2 _15588_ (.A(_06631_),
    .B(_06656_),
    .Y(_06657_));
 sky130_fd_sc_hd__a21oi_4 _15589_ (.A1(_06540_),
    .A2(_06565_),
    .B1(_06657_),
    .Y(_06658_));
 sky130_fd_sc_hd__and3_1 _15590_ (.A(_06540_),
    .B(_06565_),
    .C(_06657_),
    .X(_06660_));
 sky130_fd_sc_hd__or2_4 _15591_ (.A(_06658_),
    .B(_06660_),
    .X(_06661_));
 sky130_fd_sc_hd__a31o_1 _15592_ (.A1(net146),
    .A2(net188),
    .A3(_06557_),
    .B1(_06555_),
    .X(_06662_));
 sky130_fd_sc_hd__nand2_2 _15593_ (.A(_06562_),
    .B(_06662_),
    .Y(_06663_));
 sky130_fd_sc_hd__or2_1 _15594_ (.A(_06562_),
    .B(_06662_),
    .X(_06664_));
 sky130_fd_sc_hd__nand2_1 _15595_ (.A(_06663_),
    .B(_06664_),
    .Y(_06665_));
 sky130_fd_sc_hd__nand2_1 _15596_ (.A(net142),
    .B(net188),
    .Y(_06666_));
 sky130_fd_sc_hd__or2_4 _15597_ (.A(_06665_),
    .B(_06666_),
    .X(_06667_));
 sky130_fd_sc_hd__nand2_1 _15598_ (.A(_06665_),
    .B(_06666_),
    .Y(_06668_));
 sky130_fd_sc_hd__nand2_4 _15599_ (.A(_06667_),
    .B(_06668_),
    .Y(_06669_));
 sky130_fd_sc_hd__nor2_2 _15600_ (.A(_06661_),
    .B(_06669_),
    .Y(_06671_));
 sky130_fd_sc_hd__xor2_4 _15601_ (.A(_06661_),
    .B(_06669_),
    .X(_06672_));
 sky130_fd_sc_hd__a21oi_4 _15602_ (.A1(_06478_),
    .A2(_06566_),
    .B1(_06574_),
    .Y(_06673_));
 sky130_fd_sc_hd__nand2b_1 _15603_ (.A_N(_06673_),
    .B(_06672_),
    .Y(_06674_));
 sky130_fd_sc_hd__xnor2_4 _15604_ (.A(_06672_),
    .B(_06673_),
    .Y(_06675_));
 sky130_fd_sc_hd__a21o_2 _15605_ (.A1(_06476_),
    .A2(_06568_),
    .B1(_06571_),
    .X(_06676_));
 sky130_fd_sc_hd__nand2_1 _15606_ (.A(_06675_),
    .B(_06676_),
    .Y(_06677_));
 sky130_fd_sc_hd__xor2_2 _15607_ (.A(_06675_),
    .B(_06676_),
    .X(_06678_));
 sky130_fd_sc_hd__o21a_1 _15608_ (.A1(_06576_),
    .A2(_06580_),
    .B1(_06678_),
    .X(_06679_));
 sky130_fd_sc_hd__nor3_1 _15609_ (.A(_06576_),
    .B(_06580_),
    .C(_06678_),
    .Y(_06680_));
 sky130_fd_sc_hd__nor2_2 _15610_ (.A(_06679_),
    .B(_06680_),
    .Y(_06682_));
 sky130_fd_sc_hd__a21o_2 _15611_ (.A1(_06529_),
    .A2(_06584_),
    .B1(_06582_),
    .X(_06683_));
 sky130_fd_sc_hd__o21a_1 _15612_ (.A1(_06682_),
    .A2(_06683_),
    .B1(net281),
    .X(_06684_));
 sky130_fd_sc_hd__a21boi_4 _15613_ (.A1(_06682_),
    .A2(_06683_),
    .B1_N(_06684_),
    .Y(_06685_));
 sky130_fd_sc_hd__and2_1 _15614_ (.A(_02417_),
    .B(_02491_),
    .X(_06686_));
 sky130_fd_sc_hd__or3_4 _15615_ (.A(_02492_),
    .B(net256),
    .C(_06686_),
    .X(_06687_));
 sky130_fd_sc_hd__a21boi_1 _15616_ (.A1(net500),
    .A2(net272),
    .B1_N(net818),
    .Y(_06688_));
 sky130_fd_sc_hd__or3b_1 _15617_ (.A(net818),
    .B(net269),
    .C_N(net500),
    .X(_06689_));
 sky130_fd_sc_hd__nand2b_1 _15618_ (.A_N(_06688_),
    .B(_06689_),
    .Y(_06690_));
 sky130_fd_sc_hd__a211o_1 _15619_ (.A1(_06508_),
    .A2(_06509_),
    .B1(_06593_),
    .C1(_06506_),
    .X(_06691_));
 sky130_fd_sc_hd__and2_1 _15620_ (.A(_06595_),
    .B(_06691_),
    .X(_06693_));
 sky130_fd_sc_hd__xnor2_1 _15621_ (.A(_06690_),
    .B(_06693_),
    .Y(_06694_));
 sky130_fd_sc_hd__nand2_1 _15622_ (.A(_01065_),
    .B(_05784_),
    .Y(_06695_));
 sky130_fd_sc_hd__xor2_2 _15623_ (.A(_05809_),
    .B(_06695_),
    .X(_06696_));
 sky130_fd_sc_hd__nor2_1 _15624_ (.A(net816),
    .B(_05859_),
    .Y(_06697_));
 sky130_fd_sc_hd__a22o_1 _15625_ (.A1(_01064_),
    .A2(net237),
    .B1(net231),
    .B2(net819),
    .X(_06698_));
 sky130_fd_sc_hd__a211oi_1 _15626_ (.A1(_05784_),
    .A2(net240),
    .B1(_06698_),
    .C1(net242),
    .Y(_06699_));
 sky130_fd_sc_hd__or2_2 _15627_ (.A(net575),
    .B(_06057_),
    .X(_06700_));
 sky130_fd_sc_hd__and2_1 _15628_ (.A(net558),
    .B(_06700_),
    .X(_06701_));
 sky130_fd_sc_hd__mux4_1 _15629_ (.A0(_06059_),
    .A1(_06061_),
    .A2(_06081_),
    .A3(_06083_),
    .S0(net299),
    .S1(net303),
    .X(_06702_));
 sky130_fd_sc_hd__a21o_1 _15630_ (.A1(net309),
    .A2(_06702_),
    .B1(net241),
    .X(_06704_));
 sky130_fd_sc_hd__o32a_1 _15631_ (.A1(net249),
    .A2(_05860_),
    .A3(_06697_),
    .B1(_06701_),
    .B2(_06704_),
    .X(_06705_));
 sky130_fd_sc_hd__o311a_1 _15632_ (.A1(net558),
    .A2(net210),
    .A3(_04000_),
    .B1(_06699_),
    .C1(_06705_),
    .X(_06706_));
 sky130_fd_sc_hd__o21ai_2 _15633_ (.A1(net253),
    .A2(_06696_),
    .B1(_06706_),
    .Y(_06707_));
 sky130_fd_sc_hd__a211oi_1 _15634_ (.A1(net230),
    .A2(_06694_),
    .B1(_06707_),
    .C1(_06685_),
    .Y(_06708_));
 sky130_fd_sc_hd__a22o_1 _15635_ (.A1(net818),
    .A2(net243),
    .B1(_06687_),
    .B2(_06708_),
    .X(_06709_));
 sky130_fd_sc_hd__inv_2 _15636_ (.A(_06709_),
    .Y(_08685_));
 sky130_fd_sc_hd__a21bo_1 _15637_ (.A1(net452),
    .A2(net313),
    .B1_N(net490),
    .X(_06710_));
 sky130_fd_sc_hd__nor2_1 _15638_ (.A(net267),
    .B(_06710_),
    .Y(_06711_));
 sky130_fd_sc_hd__or2_4 _15639_ (.A(net267),
    .B(_06710_),
    .X(_06712_));
 sky130_fd_sc_hd__nand2_2 _15640_ (.A(net188),
    .B(net223),
    .Y(_06714_));
 sky130_fd_sc_hd__or2_4 _15641_ (.A(_06099_),
    .B(_06714_),
    .X(_06715_));
 sky130_fd_sc_hd__a22o_1 _15642_ (.A1(net140),
    .A2(net188),
    .B1(net224),
    .B2(net153),
    .X(_06716_));
 sky130_fd_sc_hd__nand2_2 _15643_ (.A(_06715_),
    .B(_06716_),
    .Y(_06717_));
 sky130_fd_sc_hd__a22o_1 _15644_ (.A1(net144),
    .A2(_06530_),
    .B1(net182),
    .B2(net149),
    .X(_06718_));
 sky130_fd_sc_hd__nor3_1 _15645_ (.A(_06042_),
    .B(_06533_),
    .C(net181),
    .Y(_06719_));
 sky130_fd_sc_hd__o31a_1 _15646_ (.A1(_06042_),
    .A2(_06533_),
    .A3(net181),
    .B1(_06718_),
    .X(_06720_));
 sky130_fd_sc_hd__nand2_1 _15647_ (.A(_06103_),
    .B(net131),
    .Y(_06721_));
 sky130_fd_sc_hd__xnor2_2 _15648_ (.A(_06720_),
    .B(_06721_),
    .Y(_06722_));
 sky130_fd_sc_hd__a31o_2 _15649_ (.A1(net144),
    .A2(net131),
    .A3(_06621_),
    .B1(_06620_),
    .X(_06723_));
 sky130_fd_sc_hd__and2_2 _15650_ (.A(_06722_),
    .B(_06723_),
    .X(_06725_));
 sky130_fd_sc_hd__xnor2_2 _15651_ (.A(_06722_),
    .B(_06723_),
    .Y(_06726_));
 sky130_fd_sc_hd__nor2_2 _15652_ (.A(_06717_),
    .B(_06726_),
    .Y(_06727_));
 sky130_fd_sc_hd__and2_1 _15653_ (.A(_06717_),
    .B(_06726_),
    .X(_06728_));
 sky130_fd_sc_hd__nor2_2 _15654_ (.A(_06727_),
    .B(_06728_),
    .Y(_06729_));
 sky130_fd_sc_hd__and3_1 _15655_ (.A(_06614_),
    .B(_06627_),
    .C(_06729_),
    .X(_06730_));
 sky130_fd_sc_hd__xnor2_2 _15656_ (.A(_06628_),
    .B(_06729_),
    .Y(_06731_));
 sky130_fd_sc_hd__and2_4 _15657_ (.A(net807),
    .B(_06642_),
    .X(_06732_));
 sky130_fd_sc_hd__nand2_8 _15658_ (.A(net808),
    .B(_06642_),
    .Y(_06733_));
 sky130_fd_sc_hd__nand2_2 _15659_ (.A(net154),
    .B(net174),
    .Y(_06734_));
 sky130_fd_sc_hd__and3_1 _15660_ (.A(net154),
    .B(_06389_),
    .C(net174),
    .X(_06736_));
 sky130_fd_sc_hd__xnor2_4 _15661_ (.A(_06389_),
    .B(_06734_),
    .Y(_06737_));
 sky130_fd_sc_hd__nand2_1 _15662_ (.A(net146),
    .B(net177),
    .Y(_06738_));
 sky130_fd_sc_hd__xnor2_2 _15663_ (.A(_06737_),
    .B(_06738_),
    .Y(_06739_));
 sky130_fd_sc_hd__nor2_8 _15664_ (.A(_06247_),
    .B(_06305_),
    .Y(_06740_));
 sky130_fd_sc_hd__nand2_1 _15665_ (.A(_06633_),
    .B(_06740_),
    .Y(_06741_));
 sky130_fd_sc_hd__xnor2_4 _15666_ (.A(_06633_),
    .B(_06740_),
    .Y(_06742_));
 sky130_fd_sc_hd__nand2_2 _15667_ (.A(net136),
    .B(net193),
    .Y(_06743_));
 sky130_fd_sc_hd__xor2_4 _15668_ (.A(_06742_),
    .B(_06743_),
    .X(_06744_));
 sky130_fd_sc_hd__a21bo_4 _15669_ (.A1(_06632_),
    .A2(_06636_),
    .B1_N(_06634_),
    .X(_06745_));
 sky130_fd_sc_hd__nand2_2 _15670_ (.A(_06744_),
    .B(_06745_),
    .Y(_06747_));
 sky130_fd_sc_hd__xor2_4 _15671_ (.A(_06744_),
    .B(_06745_),
    .X(_06748_));
 sky130_fd_sc_hd__nand2_2 _15672_ (.A(_06739_),
    .B(_06748_),
    .Y(_06749_));
 sky130_fd_sc_hd__xnor2_1 _15673_ (.A(_06739_),
    .B(_06748_),
    .Y(_06750_));
 sky130_fd_sc_hd__and2_2 _15674_ (.A(_06625_),
    .B(_06750_),
    .X(_06751_));
 sky130_fd_sc_hd__nor2_2 _15675_ (.A(_06625_),
    .B(_06750_),
    .Y(_06752_));
 sky130_fd_sc_hd__inv_2 _15676_ (.A(_06752_),
    .Y(_06753_));
 sky130_fd_sc_hd__a211o_2 _15677_ (.A1(_06640_),
    .A2(_06652_),
    .B1(_06751_),
    .C1(_06752_),
    .X(_06754_));
 sky130_fd_sc_hd__o211ai_4 _15678_ (.A1(_06751_),
    .A2(_06752_),
    .B1(_06640_),
    .C1(_06652_),
    .Y(_06755_));
 sky130_fd_sc_hd__and3_2 _15679_ (.A(_06731_),
    .B(_06754_),
    .C(_06755_),
    .X(_06756_));
 sky130_fd_sc_hd__a21oi_4 _15680_ (.A1(_06754_),
    .A2(_06755_),
    .B1(_06731_),
    .Y(_06758_));
 sky130_fd_sc_hd__a21oi_4 _15681_ (.A1(_06631_),
    .A2(_06656_),
    .B1(_06630_),
    .Y(_06759_));
 sky130_fd_sc_hd__nor3_4 _15682_ (.A(_06756_),
    .B(_06758_),
    .C(_06759_),
    .Y(_06760_));
 sky130_fd_sc_hd__o21a_1 _15683_ (.A1(_06756_),
    .A2(_06758_),
    .B1(_06759_),
    .X(_06761_));
 sky130_fd_sc_hd__o21ba_1 _15684_ (.A1(_06647_),
    .A2(_06650_),
    .B1_N(_06646_),
    .X(_06762_));
 sky130_fd_sc_hd__or3b_1 _15685_ (.A(_06762_),
    .B(_06653_),
    .C_N(_06654_),
    .X(_06763_));
 sky130_fd_sc_hd__xnor2_1 _15686_ (.A(_06655_),
    .B(_06762_),
    .Y(_06764_));
 sky130_fd_sc_hd__or3b_2 _15687_ (.A(_06048_),
    .B(net183),
    .C_N(_06764_),
    .X(_06765_));
 sky130_fd_sc_hd__a21o_1 _15688_ (.A1(net141),
    .A2(net184),
    .B1(_06764_),
    .X(_06766_));
 sky130_fd_sc_hd__nand2_2 _15689_ (.A(_06765_),
    .B(_06766_),
    .Y(_06767_));
 sky130_fd_sc_hd__or3_4 _15690_ (.A(_06760_),
    .B(_06761_),
    .C(_06767_),
    .X(_06769_));
 sky130_fd_sc_hd__o21ai_4 _15691_ (.A1(_06760_),
    .A2(_06761_),
    .B1(_06767_),
    .Y(_06770_));
 sky130_fd_sc_hd__o211a_2 _15692_ (.A1(_06658_),
    .A2(_06671_),
    .B1(_06769_),
    .C1(_06770_),
    .X(_06771_));
 sky130_fd_sc_hd__a211oi_4 _15693_ (.A1(_06769_),
    .A2(_06770_),
    .B1(_06658_),
    .C1(_06671_),
    .Y(_06772_));
 sky130_fd_sc_hd__a211oi_4 _15694_ (.A1(_06663_),
    .A2(_06667_),
    .B1(_06771_),
    .C1(_06772_),
    .Y(_06773_));
 sky130_fd_sc_hd__o211a_1 _15695_ (.A1(_06771_),
    .A2(_06772_),
    .B1(_06663_),
    .C1(_06667_),
    .X(_06774_));
 sky130_fd_sc_hd__a211oi_2 _15696_ (.A1(_06674_),
    .A2(_06677_),
    .B1(_06773_),
    .C1(_06774_),
    .Y(_06775_));
 sky130_fd_sc_hd__o211a_1 _15697_ (.A1(_06773_),
    .A2(_06774_),
    .B1(_06674_),
    .C1(_06677_),
    .X(_06776_));
 sky130_fd_sc_hd__nor2_1 _15698_ (.A(_06775_),
    .B(_06776_),
    .Y(_06777_));
 sky130_fd_sc_hd__a21oi_1 _15699_ (.A1(_06682_),
    .A2(_06683_),
    .B1(_06679_),
    .Y(_06778_));
 sky130_fd_sc_hd__xnor2_1 _15700_ (.A(_06777_),
    .B(_06778_),
    .Y(_06780_));
 sky130_fd_sc_hd__a21o_1 _15701_ (.A1(_02381_),
    .A2(_02494_),
    .B1(_02493_),
    .X(_06781_));
 sky130_fd_sc_hd__a21o_1 _15702_ (.A1(net490),
    .A2(net272),
    .B1(_03269_),
    .X(_06782_));
 sky130_fd_sc_hd__or3b_4 _15703_ (.A(net808),
    .B(net270),
    .C_N(net490),
    .X(_06783_));
 sky130_fd_sc_hd__a31o_2 _15704_ (.A1(_06595_),
    .A2(_06689_),
    .A3(_06691_),
    .B1(_06688_),
    .X(_06784_));
 sky130_fd_sc_hd__nand3_1 _15705_ (.A(_06782_),
    .B(_06783_),
    .C(_06784_),
    .Y(_06785_));
 sky130_fd_sc_hd__a21o_1 _15706_ (.A1(_06782_),
    .A2(_06783_),
    .B1(_06784_),
    .X(_06786_));
 sky130_fd_sc_hd__nand3_1 _15707_ (.A(_00937_),
    .B(_05783_),
    .C(_05810_),
    .Y(_06787_));
 sky130_fd_sc_hd__a21o_1 _15708_ (.A1(_00937_),
    .A2(_05783_),
    .B1(_05810_),
    .X(_06788_));
 sky130_fd_sc_hd__nor2_1 _15709_ (.A(net807),
    .B(_05860_),
    .Y(_06789_));
 sky130_fd_sc_hd__or3_1 _15710_ (.A(net249),
    .B(_05861_),
    .C(_06789_),
    .X(_06791_));
 sky130_fd_sc_hd__nor2_1 _15711_ (.A(net577),
    .B(_06157_),
    .Y(_06792_));
 sky130_fd_sc_hd__a211o_1 _15712_ (.A1(net577),
    .A2(_06131_),
    .B1(_06792_),
    .C1(net203),
    .X(_06793_));
 sky130_fd_sc_hd__a221o_1 _15713_ (.A1(_05783_),
    .A2(net240),
    .B1(net231),
    .B2(net807),
    .C1(net242),
    .X(_06794_));
 sky130_fd_sc_hd__a21oi_1 _15714_ (.A1(_00936_),
    .A2(net237),
    .B1(_06794_),
    .Y(_06795_));
 sky130_fd_sc_hd__or2_2 _15715_ (.A(net575),
    .B(_06125_),
    .X(_06796_));
 sky130_fd_sc_hd__o2111a_1 _15716_ (.A1(_05980_),
    .A2(_06796_),
    .B1(_06795_),
    .C1(_06793_),
    .D1(_06791_),
    .X(_06797_));
 sky130_fd_sc_hd__o31ai_1 _15717_ (.A1(net544),
    .A2(net207),
    .A3(_04143_),
    .B1(_06797_),
    .Y(_06798_));
 sky130_fd_sc_hd__a31o_1 _15718_ (.A1(net254),
    .A2(_06787_),
    .A3(_06788_),
    .B1(_06798_),
    .X(_06799_));
 sky130_fd_sc_hd__a31o_2 _15719_ (.A1(net230),
    .A2(_06785_),
    .A3(_06786_),
    .B1(_06799_),
    .X(_06800_));
 sky130_fd_sc_hd__a31o_1 _15720_ (.A1(_02495_),
    .A2(net261),
    .A3(_06781_),
    .B1(_06800_),
    .X(_06802_));
 sky130_fd_sc_hd__a21o_2 _15721_ (.A1(net281),
    .A2(_06780_),
    .B1(_06802_),
    .X(_06803_));
 sky130_fd_sc_hd__o21a_1 _15722_ (.A1(_03269_),
    .A2(_05880_),
    .B1(_06803_),
    .X(_08686_));
 sky130_fd_sc_hd__nor2_4 _15723_ (.A(net139),
    .B(_06553_),
    .Y(_06804_));
 sky130_fd_sc_hd__and2_2 _15724_ (.A(net478),
    .B(net226),
    .X(_06805_));
 sky130_fd_sc_hd__nand2_2 _15725_ (.A(net478),
    .B(net225),
    .Y(_06806_));
 sky130_fd_sc_hd__and4_4 _15726_ (.A(net153),
    .B(net149),
    .C(net224),
    .D(net172),
    .X(_06807_));
 sky130_fd_sc_hd__o22a_2 _15727_ (.A1(_05987_),
    .A2(_06712_),
    .B1(_06806_),
    .B2(_05920_),
    .X(_06808_));
 sky130_fd_sc_hd__nor2_4 _15728_ (.A(_06807_),
    .B(_06808_),
    .Y(_06809_));
 sky130_fd_sc_hd__nand2_4 _15729_ (.A(_06804_),
    .B(_06809_),
    .Y(_06810_));
 sky130_fd_sc_hd__xnor2_4 _15730_ (.A(_06804_),
    .B(_06809_),
    .Y(_06812_));
 sky130_fd_sc_hd__or2_1 _15731_ (.A(_06715_),
    .B(_06812_),
    .X(_06813_));
 sky130_fd_sc_hd__xnor2_4 _15732_ (.A(_06715_),
    .B(_06812_),
    .Y(_06814_));
 sky130_fd_sc_hd__a22o_1 _15733_ (.A1(_06103_),
    .A2(_06530_),
    .B1(net182),
    .B2(net143),
    .X(_06815_));
 sky130_fd_sc_hd__or4_4 _15734_ (.A(_06042_),
    .B(net138),
    .C(net186),
    .D(net181),
    .X(_06816_));
 sky130_fd_sc_hd__nand2_4 _15735_ (.A(_06815_),
    .B(_06816_),
    .Y(_06817_));
 sky130_fd_sc_hd__nand2_4 _15736_ (.A(net199),
    .B(net131),
    .Y(_06818_));
 sky130_fd_sc_hd__xnor2_4 _15737_ (.A(_06817_),
    .B(_06818_),
    .Y(_06819_));
 sky130_fd_sc_hd__a31o_4 _15738_ (.A1(_06103_),
    .A2(net131),
    .A3(_06718_),
    .B1(_06719_),
    .X(_06820_));
 sky130_fd_sc_hd__and2b_4 _15739_ (.A_N(_06819_),
    .B(_06820_),
    .X(_06821_));
 sky130_fd_sc_hd__xor2_4 _15740_ (.A(_06819_),
    .B(_06820_),
    .X(_06823_));
 sky130_fd_sc_hd__xnor2_4 _15741_ (.A(_06814_),
    .B(_06823_),
    .Y(_06824_));
 sky130_fd_sc_hd__nor3_1 _15742_ (.A(_06717_),
    .B(_06726_),
    .C(_06824_),
    .Y(_06825_));
 sky130_fd_sc_hd__xor2_2 _15743_ (.A(_06727_),
    .B(_06824_),
    .X(_06826_));
 sky130_fd_sc_hd__and2_4 _15744_ (.A(net797),
    .B(net227),
    .X(_06827_));
 sky130_fd_sc_hd__nand2_8 _15745_ (.A(net797),
    .B(net225),
    .Y(_06828_));
 sky130_fd_sc_hd__or2_4 _15746_ (.A(net201),
    .B(_06828_),
    .X(_06829_));
 sky130_fd_sc_hd__a2bb2o_1 _15747_ (.A1_N(net201),
    .A2_N(_06465_),
    .B1(_06827_),
    .B2(net155),
    .X(_06830_));
 sky130_fd_sc_hd__o21a_2 _15748_ (.A1(_06467_),
    .A2(_06829_),
    .B1(_06830_),
    .X(_06831_));
 sky130_fd_sc_hd__nand2_2 _15749_ (.A(net147),
    .B(net174),
    .Y(_06832_));
 sky130_fd_sc_hd__and3_1 _15750_ (.A(_05990_),
    .B(_06732_),
    .C(_06831_),
    .X(_06834_));
 sky130_fd_sc_hd__xor2_4 _15751_ (.A(_06831_),
    .B(_06832_),
    .X(_06835_));
 sky130_fd_sc_hd__nor2_8 _15752_ (.A(net191),
    .B(net189),
    .Y(_06836_));
 sky130_fd_sc_hd__o22a_1 _15753_ (.A1(_06305_),
    .A2(net192),
    .B1(net190),
    .B2(net196),
    .X(_06837_));
 sky130_fd_sc_hd__a21oi_4 _15754_ (.A1(_06740_),
    .A2(_06836_),
    .B1(_06837_),
    .Y(_06838_));
 sky130_fd_sc_hd__nor2_4 _15755_ (.A(_06236_),
    .B(net133),
    .Y(_06839_));
 sky130_fd_sc_hd__xnor2_4 _15756_ (.A(_06838_),
    .B(_06839_),
    .Y(_06840_));
 sky130_fd_sc_hd__o21a_2 _15757_ (.A1(_06742_),
    .A2(_06743_),
    .B1(_06741_),
    .X(_06841_));
 sky130_fd_sc_hd__or2_2 _15758_ (.A(_06840_),
    .B(_06841_),
    .X(_06842_));
 sky130_fd_sc_hd__xnor2_4 _15759_ (.A(_06840_),
    .B(_06841_),
    .Y(_06843_));
 sky130_fd_sc_hd__xor2_4 _15760_ (.A(_06835_),
    .B(_06843_),
    .X(_06845_));
 sky130_fd_sc_hd__and2_1 _15761_ (.A(_06725_),
    .B(_06845_),
    .X(_06846_));
 sky130_fd_sc_hd__xnor2_2 _15762_ (.A(_06725_),
    .B(_06845_),
    .Y(_06847_));
 sky130_fd_sc_hd__a21oi_4 _15763_ (.A1(_06747_),
    .A2(_06749_),
    .B1(_06847_),
    .Y(_06848_));
 sky130_fd_sc_hd__and3_1 _15764_ (.A(_06747_),
    .B(_06749_),
    .C(_06847_),
    .X(_06849_));
 sky130_fd_sc_hd__nor3_2 _15765_ (.A(_06826_),
    .B(_06848_),
    .C(_06849_),
    .Y(_06850_));
 sky130_fd_sc_hd__o21a_1 _15766_ (.A1(_06848_),
    .A2(_06849_),
    .B1(_06826_),
    .X(_06851_));
 sky130_fd_sc_hd__nor2_1 _15767_ (.A(_06850_),
    .B(_06851_),
    .Y(_06852_));
 sky130_fd_sc_hd__o21a_1 _15768_ (.A1(_06730_),
    .A2(_06756_),
    .B1(_06852_),
    .X(_06853_));
 sky130_fd_sc_hd__nor3_1 _15769_ (.A(_06730_),
    .B(_06756_),
    .C(_06852_),
    .Y(_06854_));
 sky130_fd_sc_hd__a31oi_2 _15770_ (.A1(net146),
    .A2(net178),
    .A3(_06737_),
    .B1(_06736_),
    .Y(_06856_));
 sky130_fd_sc_hd__a21oi_1 _15771_ (.A1(_06753_),
    .A2(_06754_),
    .B1(_06856_),
    .Y(_06857_));
 sky130_fd_sc_hd__and3_1 _15772_ (.A(_06753_),
    .B(_06754_),
    .C(_06856_),
    .X(_06858_));
 sky130_fd_sc_hd__nor2_1 _15773_ (.A(_06857_),
    .B(_06858_),
    .Y(_06859_));
 sky130_fd_sc_hd__nand2_1 _15774_ (.A(net142),
    .B(net178),
    .Y(_06860_));
 sky130_fd_sc_hd__xor2_1 _15775_ (.A(_06859_),
    .B(_06860_),
    .X(_06861_));
 sky130_fd_sc_hd__nor3_1 _15776_ (.A(_06853_),
    .B(_06854_),
    .C(_06861_),
    .Y(_06862_));
 sky130_fd_sc_hd__o21a_1 _15777_ (.A1(_06853_),
    .A2(_06854_),
    .B1(_06861_),
    .X(_06863_));
 sky130_fd_sc_hd__or2_1 _15778_ (.A(_06862_),
    .B(_06863_),
    .X(_06864_));
 sky130_fd_sc_hd__nand2b_1 _15779_ (.A_N(_06760_),
    .B(_06769_),
    .Y(_06865_));
 sky130_fd_sc_hd__and2b_1 _15780_ (.A_N(_06864_),
    .B(_06865_),
    .X(_06867_));
 sky130_fd_sc_hd__xnor2_1 _15781_ (.A(_06864_),
    .B(_06865_),
    .Y(_06868_));
 sky130_fd_sc_hd__nand2_1 _15782_ (.A(_06763_),
    .B(_06765_),
    .Y(_06869_));
 sky130_fd_sc_hd__and2_2 _15783_ (.A(_06868_),
    .B(_06869_),
    .X(_06870_));
 sky130_fd_sc_hd__nor2_1 _15784_ (.A(_06868_),
    .B(_06869_),
    .Y(_06871_));
 sky130_fd_sc_hd__or2_4 _15785_ (.A(_06870_),
    .B(_06871_),
    .X(_06872_));
 sky130_fd_sc_hd__or2_4 _15786_ (.A(_06771_),
    .B(_06773_),
    .X(_06873_));
 sky130_fd_sc_hd__or3b_1 _15787_ (.A(_06870_),
    .B(_06871_),
    .C_N(_06873_),
    .X(_06874_));
 sky130_fd_sc_hd__xnor2_4 _15788_ (.A(_06872_),
    .B(_06873_),
    .Y(_06875_));
 sky130_fd_sc_hd__o21ba_1 _15789_ (.A1(_06679_),
    .A2(_06775_),
    .B1_N(_06776_),
    .X(_06876_));
 sky130_fd_sc_hd__a31o_2 _15790_ (.A1(_06682_),
    .A2(_06683_),
    .A3(_06777_),
    .B1(_06876_),
    .X(_06878_));
 sky130_fd_sc_hd__o21ai_1 _15791_ (.A1(_06875_),
    .A2(_06878_),
    .B1(net281),
    .Y(_06879_));
 sky130_fd_sc_hd__a21o_2 _15792_ (.A1(_06875_),
    .A2(_06878_),
    .B1(_06879_),
    .X(_06880_));
 sky130_fd_sc_hd__nor2_1 _15793_ (.A(_02344_),
    .B(_02496_),
    .Y(_06881_));
 sky130_fd_sc_hd__or3b_4 _15794_ (.A(net256),
    .B(_06881_),
    .C_N(_02497_),
    .X(_06882_));
 sky130_fd_sc_hd__a21bo_1 _15795_ (.A1(net478),
    .A2(net276),
    .B1_N(net796),
    .X(_06883_));
 sky130_fd_sc_hd__or3b_1 _15796_ (.A(net798),
    .B(net270),
    .C_N(net478),
    .X(_06884_));
 sky130_fd_sc_hd__nand2_1 _15797_ (.A(_06883_),
    .B(_06884_),
    .Y(_06885_));
 sky130_fd_sc_hd__a21boi_4 _15798_ (.A1(_06783_),
    .A2(_06784_),
    .B1_N(_06782_),
    .Y(_06886_));
 sky130_fd_sc_hd__a21oi_1 _15799_ (.A1(_06885_),
    .A2(_06886_),
    .B1(net229),
    .Y(_06887_));
 sky130_fd_sc_hd__o21ai_1 _15800_ (.A1(_06885_),
    .A2(_06886_),
    .B1(_06887_),
    .Y(_06889_));
 sky130_fd_sc_hd__and2_1 _15801_ (.A(_00654_),
    .B(_05782_),
    .X(_06890_));
 sky130_fd_sc_hd__xnor2_1 _15802_ (.A(_05811_),
    .B(_06890_),
    .Y(_06891_));
 sky130_fd_sc_hd__a221o_1 _15803_ (.A1(_05782_),
    .A2(net239),
    .B1(net234),
    .B2(net796),
    .C1(net243),
    .X(_06892_));
 sky130_fd_sc_hd__a21oi_1 _15804_ (.A1(_00653_),
    .A2(net236),
    .B1(_06892_),
    .Y(_06893_));
 sky130_fd_sc_hd__nor2_1 _15805_ (.A(net576),
    .B(_06227_),
    .Y(_06894_));
 sky130_fd_sc_hd__o21ai_1 _15806_ (.A1(net301),
    .A2(_06213_),
    .B1(net308),
    .Y(_06895_));
 sky130_fd_sc_hd__o21a_1 _15807_ (.A1(net575),
    .A2(_06215_),
    .B1(net559),
    .X(_06896_));
 sky130_fd_sc_hd__nor2_1 _15808_ (.A(net241),
    .B(_06896_),
    .Y(_06897_));
 sky130_fd_sc_hd__o21ai_1 _15809_ (.A1(_06894_),
    .A2(_06895_),
    .B1(_06897_),
    .Y(_06898_));
 sky130_fd_sc_hd__o311a_1 _15810_ (.A1(net544),
    .A2(net207),
    .A3(_04271_),
    .B1(_06893_),
    .C1(_06898_),
    .X(_06900_));
 sky130_fd_sc_hd__nor2_1 _15811_ (.A(net796),
    .B(_05861_),
    .Y(_06901_));
 sky130_fd_sc_hd__o31a_1 _15812_ (.A1(net251),
    .A2(_05862_),
    .A3(_06901_),
    .B1(_06900_),
    .X(_06902_));
 sky130_fd_sc_hd__o211a_1 _15813_ (.A1(_05841_),
    .A2(_06891_),
    .B1(_06902_),
    .C1(_06889_),
    .X(_06903_));
 sky130_fd_sc_hd__a32o_1 _15814_ (.A1(_06880_),
    .A2(_06882_),
    .A3(_06903_),
    .B1(net243),
    .B2(net796),
    .X(_06904_));
 sky130_fd_sc_hd__clkinv_2 _15815_ (.A(_06904_),
    .Y(_08687_));
 sky130_fd_sc_hd__nor2_4 _15816_ (.A(net139),
    .B(net176),
    .Y(_06905_));
 sky130_fd_sc_hd__and2_2 _15817_ (.A(net471),
    .B(net226),
    .X(_06906_));
 sky130_fd_sc_hd__nand2_2 _15818_ (.A(net471),
    .B(net225),
    .Y(_06907_));
 sky130_fd_sc_hd__a22o_1 _15819_ (.A1(net149),
    .A2(net172),
    .B1(net170),
    .B2(_05919_),
    .X(_06908_));
 sky130_fd_sc_hd__or4_1 _15820_ (.A(_05920_),
    .B(_05987_),
    .C(_06806_),
    .D(net169),
    .X(_06910_));
 sky130_fd_sc_hd__and4_1 _15821_ (.A(net143),
    .B(net224),
    .C(_06908_),
    .D(_06910_),
    .X(_06911_));
 sky130_fd_sc_hd__a22o_1 _15822_ (.A1(net143),
    .A2(net224),
    .B1(_06908_),
    .B2(_06910_),
    .X(_06912_));
 sky130_fd_sc_hd__and2b_4 _15823_ (.A_N(_06911_),
    .B(_06912_),
    .X(_06913_));
 sky130_fd_sc_hd__nand2_1 _15824_ (.A(_06905_),
    .B(_06913_),
    .Y(_06914_));
 sky130_fd_sc_hd__xnor2_4 _15825_ (.A(_06905_),
    .B(_06913_),
    .Y(_06915_));
 sky130_fd_sc_hd__nor2_1 _15826_ (.A(_06810_),
    .B(_06915_),
    .Y(_06916_));
 sky130_fd_sc_hd__xor2_4 _15827_ (.A(_06810_),
    .B(_06915_),
    .X(_06917_));
 sky130_fd_sc_hd__o21ai_4 _15828_ (.A1(_06817_),
    .A2(_06818_),
    .B1(_06816_),
    .Y(_06918_));
 sky130_fd_sc_hd__o22a_1 _15829_ (.A1(_06184_),
    .A2(net186),
    .B1(net180),
    .B2(_06104_),
    .X(_06919_));
 sky130_fd_sc_hd__or4_1 _15830_ (.A(net138),
    .B(_06184_),
    .C(net185),
    .D(net180),
    .X(_06921_));
 sky130_fd_sc_hd__and2b_2 _15831_ (.A_N(_06919_),
    .B(_06921_),
    .X(_06922_));
 sky130_fd_sc_hd__xnor2_4 _15832_ (.A(_06449_),
    .B(_06922_),
    .Y(_06923_));
 sky130_fd_sc_hd__nand2_1 _15833_ (.A(_06807_),
    .B(_06923_),
    .Y(_06924_));
 sky130_fd_sc_hd__xnor2_4 _15834_ (.A(_06807_),
    .B(_06923_),
    .Y(_06925_));
 sky130_fd_sc_hd__nand2b_1 _15835_ (.A_N(_06925_),
    .B(_06918_),
    .Y(_06926_));
 sky130_fd_sc_hd__xnor2_4 _15836_ (.A(_06918_),
    .B(_06925_),
    .Y(_06927_));
 sky130_fd_sc_hd__xnor2_2 _15837_ (.A(_06917_),
    .B(_06927_),
    .Y(_06928_));
 sky130_fd_sc_hd__o21a_2 _15838_ (.A1(_06814_),
    .A2(_06823_),
    .B1(_06813_),
    .X(_06929_));
 sky130_fd_sc_hd__nor2_1 _15839_ (.A(_06928_),
    .B(_06929_),
    .Y(_06930_));
 sky130_fd_sc_hd__nand2_1 _15840_ (.A(_06928_),
    .B(_06929_),
    .Y(_06932_));
 sky130_fd_sc_hd__xnor2_1 _15841_ (.A(_06928_),
    .B(_06929_),
    .Y(_06933_));
 sky130_fd_sc_hd__o21ai_4 _15842_ (.A1(_06835_),
    .A2(_06843_),
    .B1(_06842_),
    .Y(_06934_));
 sky130_fd_sc_hd__and2_4 _15843_ (.A(net784),
    .B(net225),
    .X(_06935_));
 sky130_fd_sc_hd__nand2_4 _15844_ (.A(net784),
    .B(net225),
    .Y(_06936_));
 sky130_fd_sc_hd__or2_1 _15845_ (.A(net200),
    .B(_06936_),
    .X(_06937_));
 sky130_fd_sc_hd__and3_2 _15846_ (.A(net155),
    .B(_06554_),
    .C(_06935_),
    .X(_06938_));
 sky130_fd_sc_hd__a21oi_2 _15847_ (.A1(net155),
    .A2(_06935_),
    .B1(_06554_),
    .Y(_06939_));
 sky130_fd_sc_hd__nor2_4 _15848_ (.A(_06938_),
    .B(_06939_),
    .Y(_06940_));
 sky130_fd_sc_hd__nand2_2 _15849_ (.A(net147),
    .B(_06827_),
    .Y(_06941_));
 sky130_fd_sc_hd__xor2_4 _15850_ (.A(_06940_),
    .B(_06941_),
    .X(_06943_));
 sky130_fd_sc_hd__nor2_8 _15851_ (.A(_06305_),
    .B(net134),
    .Y(_06944_));
 sky130_fd_sc_hd__nand2_1 _15852_ (.A(_06836_),
    .B(_06944_),
    .Y(_06945_));
 sky130_fd_sc_hd__xnor2_4 _15853_ (.A(_06836_),
    .B(_06944_),
    .Y(_06946_));
 sky130_fd_sc_hd__nand2_4 _15854_ (.A(net136),
    .B(net188),
    .Y(_06947_));
 sky130_fd_sc_hd__xnor2_4 _15855_ (.A(_06946_),
    .B(_06947_),
    .Y(_06948_));
 sky130_fd_sc_hd__a22oi_4 _15856_ (.A1(_06740_),
    .A2(_06836_),
    .B1(_06838_),
    .B2(_06839_),
    .Y(_06949_));
 sky130_fd_sc_hd__or2_1 _15857_ (.A(_06948_),
    .B(_06949_),
    .X(_06950_));
 sky130_fd_sc_hd__xnor2_4 _15858_ (.A(_06948_),
    .B(_06949_),
    .Y(_06951_));
 sky130_fd_sc_hd__xor2_4 _15859_ (.A(_06943_),
    .B(_06951_),
    .X(_06952_));
 sky130_fd_sc_hd__and2_1 _15860_ (.A(_06821_),
    .B(_06952_),
    .X(_06954_));
 sky130_fd_sc_hd__xnor2_4 _15861_ (.A(_06821_),
    .B(_06952_),
    .Y(_06955_));
 sky130_fd_sc_hd__and2b_1 _15862_ (.A_N(_06955_),
    .B(_06934_),
    .X(_06956_));
 sky130_fd_sc_hd__xnor2_4 _15863_ (.A(_06934_),
    .B(_06955_),
    .Y(_06957_));
 sky130_fd_sc_hd__xnor2_1 _15864_ (.A(_06933_),
    .B(_06957_),
    .Y(_06958_));
 sky130_fd_sc_hd__o21ai_1 _15865_ (.A1(_06825_),
    .A2(_06850_),
    .B1(_06958_),
    .Y(_06959_));
 sky130_fd_sc_hd__or3_1 _15866_ (.A(_06825_),
    .B(_06850_),
    .C(_06958_),
    .X(_06960_));
 sky130_fd_sc_hd__and2_1 _15867_ (.A(_06959_),
    .B(_06960_),
    .X(_06961_));
 sky130_fd_sc_hd__or2_1 _15868_ (.A(_06846_),
    .B(_06848_),
    .X(_06962_));
 sky130_fd_sc_hd__o21ba_1 _15869_ (.A1(_06467_),
    .A2(_06829_),
    .B1_N(_06834_),
    .X(_06963_));
 sky130_fd_sc_hd__o21ba_1 _15870_ (.A1(_06846_),
    .A2(_06848_),
    .B1_N(_06963_),
    .X(_06965_));
 sky130_fd_sc_hd__xnor2_1 _15871_ (.A(_06962_),
    .B(_06963_),
    .Y(_06966_));
 sky130_fd_sc_hd__and3_1 _15872_ (.A(net142),
    .B(net174),
    .C(_06966_),
    .X(_06967_));
 sky130_fd_sc_hd__a21oi_1 _15873_ (.A1(_06047_),
    .A2(net174),
    .B1(_06966_),
    .Y(_06968_));
 sky130_fd_sc_hd__nor2_1 _15874_ (.A(_06967_),
    .B(_06968_),
    .Y(_06969_));
 sky130_fd_sc_hd__xnor2_1 _15875_ (.A(_06961_),
    .B(_06969_),
    .Y(_06970_));
 sky130_fd_sc_hd__o21ba_1 _15876_ (.A1(_06853_),
    .A2(_06862_),
    .B1_N(_06970_),
    .X(_06971_));
 sky130_fd_sc_hd__or3b_1 _15877_ (.A(_06853_),
    .B(_06862_),
    .C_N(_06970_),
    .X(_06972_));
 sky130_fd_sc_hd__nand2b_1 _15878_ (.A_N(_06971_),
    .B(_06972_),
    .Y(_06973_));
 sky130_fd_sc_hd__o21ba_1 _15879_ (.A1(_06858_),
    .A2(_06860_),
    .B1_N(_06857_),
    .X(_06974_));
 sky130_fd_sc_hd__nor2_1 _15880_ (.A(_06973_),
    .B(_06974_),
    .Y(_06976_));
 sky130_fd_sc_hd__xnor2_1 _15881_ (.A(_06973_),
    .B(_06974_),
    .Y(_06977_));
 sky130_fd_sc_hd__o21bai_4 _15882_ (.A1(_06867_),
    .A2(_06870_),
    .B1_N(_06977_),
    .Y(_06978_));
 sky130_fd_sc_hd__or3b_2 _15883_ (.A(_06867_),
    .B(_06870_),
    .C_N(_06977_),
    .X(_06979_));
 sky130_fd_sc_hd__nand2_4 _15884_ (.A(_06978_),
    .B(_06979_),
    .Y(_06980_));
 sky130_fd_sc_hd__a21boi_4 _15885_ (.A1(_06875_),
    .A2(_06878_),
    .B1_N(_06874_),
    .Y(_06981_));
 sky130_fd_sc_hd__a21oi_2 _15886_ (.A1(_06980_),
    .A2(_06981_),
    .B1(net279),
    .Y(_06982_));
 sky130_fd_sc_hd__o21ai_4 _15887_ (.A1(_06980_),
    .A2(_06981_),
    .B1(_06982_),
    .Y(_06983_));
 sky130_fd_sc_hd__nand2_2 _15888_ (.A(_02342_),
    .B(_02497_),
    .Y(_06984_));
 sky130_fd_sc_hd__xnor2_4 _15889_ (.A(_02499_),
    .B(_06984_),
    .Y(_06985_));
 sky130_fd_sc_hd__a21bo_1 _15890_ (.A1(net471),
    .A2(net276),
    .B1_N(net785),
    .X(_06987_));
 sky130_fd_sc_hd__or3b_2 _15891_ (.A(net785),
    .B(net270),
    .C_N(net471),
    .X(_06988_));
 sky130_fd_sc_hd__o21ai_2 _15892_ (.A1(_06885_),
    .A2(_06886_),
    .B1(_06883_),
    .Y(_06989_));
 sky130_fd_sc_hd__a21oi_1 _15893_ (.A1(_06987_),
    .A2(_06988_),
    .B1(_06989_),
    .Y(_06990_));
 sky130_fd_sc_hd__a311o_1 _15894_ (.A1(_06987_),
    .A2(_06988_),
    .A3(_06989_),
    .B1(_06990_),
    .C1(net228),
    .X(_06991_));
 sky130_fd_sc_hd__and3_1 _15895_ (.A(_00220_),
    .B(_05781_),
    .C(_05813_),
    .X(_06992_));
 sky130_fd_sc_hd__a21oi_1 _15896_ (.A1(_00220_),
    .A2(_05781_),
    .B1(_05813_),
    .Y(_06993_));
 sky130_fd_sc_hd__or3_1 _15897_ (.A(net253),
    .B(_06992_),
    .C(_06993_),
    .X(_06994_));
 sky130_fd_sc_hd__nor2_1 _15898_ (.A(net786),
    .B(_05862_),
    .Y(_06995_));
 sky130_fd_sc_hd__a221o_1 _15899_ (.A1(_05781_),
    .A2(net239),
    .B1(net234),
    .B2(net786),
    .C1(net243),
    .X(_06996_));
 sky130_fd_sc_hd__a21oi_1 _15900_ (.A1(_00219_),
    .A2(net237),
    .B1(_06996_),
    .Y(_06998_));
 sky130_fd_sc_hd__mux2_1 _15901_ (.A0(_06285_),
    .A1(_06294_),
    .S(net301),
    .X(_06999_));
 sky130_fd_sc_hd__o21a_1 _15902_ (.A1(net568),
    .A2(_06293_),
    .B1(net553),
    .X(_07000_));
 sky130_fd_sc_hd__a211o_1 _15903_ (.A1(net308),
    .A2(_06999_),
    .B1(_07000_),
    .C1(net241),
    .X(_07001_));
 sky130_fd_sc_hd__o311a_1 _15904_ (.A1(net544),
    .A2(net207),
    .A3(_04408_),
    .B1(_06998_),
    .C1(_07001_),
    .X(_07002_));
 sky130_fd_sc_hd__o311a_1 _15905_ (.A1(net250),
    .A2(_05863_),
    .A3(_06995_),
    .B1(_07002_),
    .C1(_06994_),
    .X(_07003_));
 sky130_fd_sc_hd__o211a_1 _15906_ (.A1(net256),
    .A2(_06985_),
    .B1(_06991_),
    .C1(_07003_),
    .X(_07004_));
 sky130_fd_sc_hd__a22o_1 _15907_ (.A1(net785),
    .A2(net247),
    .B1(_06983_),
    .B2(_07004_),
    .X(_07005_));
 sky130_fd_sc_hd__inv_2 _15908_ (.A(_07005_),
    .Y(_08688_));
 sky130_fd_sc_hd__o21ai_4 _15909_ (.A1(_06980_),
    .A2(_06981_),
    .B1(_06978_),
    .Y(_07006_));
 sky130_fd_sc_hd__and2_2 _15910_ (.A(net461),
    .B(net225),
    .X(_07008_));
 sky130_fd_sc_hd__nand2_8 _15911_ (.A(net462),
    .B(net225),
    .Y(_07009_));
 sky130_fd_sc_hd__nand2_4 _15912_ (.A(net173),
    .B(_07008_),
    .Y(_07010_));
 sky130_fd_sc_hd__nor2_4 _15913_ (.A(_06099_),
    .B(_07010_),
    .Y(_07011_));
 sky130_fd_sc_hd__o22a_1 _15914_ (.A1(net139),
    .A2(_06733_),
    .B1(_07009_),
    .B2(_05920_),
    .X(_07012_));
 sky130_fd_sc_hd__or2_2 _15915_ (.A(_07011_),
    .B(_07012_),
    .X(_07013_));
 sky130_fd_sc_hd__a22o_1 _15916_ (.A1(net143),
    .A2(net172),
    .B1(net170),
    .B2(net148),
    .X(_07014_));
 sky130_fd_sc_hd__nand2_1 _15917_ (.A(net143),
    .B(net170),
    .Y(_07015_));
 sky130_fd_sc_hd__and4_1 _15918_ (.A(net149),
    .B(net143),
    .C(net172),
    .D(net170),
    .X(_07016_));
 sky130_fd_sc_hd__o31a_4 _15919_ (.A1(_05987_),
    .A2(net171),
    .A3(_07015_),
    .B1(_07014_),
    .X(_07017_));
 sky130_fd_sc_hd__nor2_2 _15920_ (.A(net138),
    .B(_06712_),
    .Y(_07019_));
 sky130_fd_sc_hd__xnor2_4 _15921_ (.A(_07017_),
    .B(_07019_),
    .Y(_07020_));
 sky130_fd_sc_hd__nor2_4 _15922_ (.A(_07013_),
    .B(_07020_),
    .Y(_07021_));
 sky130_fd_sc_hd__and2_1 _15923_ (.A(_07013_),
    .B(_07020_),
    .X(_07022_));
 sky130_fd_sc_hd__or2_1 _15924_ (.A(_07021_),
    .B(_07022_),
    .X(_07023_));
 sky130_fd_sc_hd__nor2_1 _15925_ (.A(_06914_),
    .B(_07023_),
    .Y(_07024_));
 sky130_fd_sc_hd__nand2_1 _15926_ (.A(_06914_),
    .B(_07023_),
    .Y(_07025_));
 sky130_fd_sc_hd__and2b_2 _15927_ (.A_N(_07024_),
    .B(_07025_),
    .X(_07026_));
 sky130_fd_sc_hd__o21ai_1 _15928_ (.A1(_06449_),
    .A2(_06919_),
    .B1(_06921_),
    .Y(_07027_));
 sky130_fd_sc_hd__a41o_1 _15929_ (.A1(_05919_),
    .A2(net149),
    .A3(_06805_),
    .A4(net170),
    .B1(_06911_),
    .X(_07028_));
 sky130_fd_sc_hd__a22o_1 _15930_ (.A1(net197),
    .A2(_06530_),
    .B1(_06617_),
    .B2(net199),
    .X(_07030_));
 sky130_fd_sc_hd__nor2_1 _15931_ (.A(net196),
    .B(net179),
    .Y(_07031_));
 sky130_fd_sc_hd__or4_1 _15932_ (.A(_06184_),
    .B(net196),
    .C(net186),
    .D(net180),
    .X(_07032_));
 sky130_fd_sc_hd__nand2_1 _15933_ (.A(_07030_),
    .B(_07032_),
    .Y(_07033_));
 sky130_fd_sc_hd__nor2_1 _15934_ (.A(net191),
    .B(_06448_),
    .Y(_07034_));
 sky130_fd_sc_hd__xnor2_1 _15935_ (.A(_07033_),
    .B(_07034_),
    .Y(_07035_));
 sky130_fd_sc_hd__and2_1 _15936_ (.A(_07028_),
    .B(_07035_),
    .X(_07036_));
 sky130_fd_sc_hd__xor2_1 _15937_ (.A(_07028_),
    .B(_07035_),
    .X(_07037_));
 sky130_fd_sc_hd__and2_2 _15938_ (.A(_07027_),
    .B(_07037_),
    .X(_07038_));
 sky130_fd_sc_hd__nor2_1 _15939_ (.A(_07027_),
    .B(_07037_),
    .Y(_07039_));
 sky130_fd_sc_hd__nor2_4 _15940_ (.A(_07038_),
    .B(_07039_),
    .Y(_07041_));
 sky130_fd_sc_hd__xnor2_4 _15941_ (.A(_07026_),
    .B(_07041_),
    .Y(_07042_));
 sky130_fd_sc_hd__a21oi_4 _15942_ (.A1(_06917_),
    .A2(_06927_),
    .B1(_06916_),
    .Y(_07043_));
 sky130_fd_sc_hd__nor2_2 _15943_ (.A(_07042_),
    .B(_07043_),
    .Y(_07044_));
 sky130_fd_sc_hd__xnor2_2 _15944_ (.A(_07042_),
    .B(_07043_),
    .Y(_07045_));
 sky130_fd_sc_hd__o21ai_1 _15945_ (.A1(_06943_),
    .A2(_06951_),
    .B1(_06950_),
    .Y(_07046_));
 sky130_fd_sc_hd__and2_4 _15946_ (.A(net776),
    .B(net226),
    .X(_07047_));
 sky130_fd_sc_hd__nand2_4 _15947_ (.A(net774),
    .B(net225),
    .Y(_07048_));
 sky130_fd_sc_hd__or2_4 _15948_ (.A(net201),
    .B(_07048_),
    .X(_07049_));
 sky130_fd_sc_hd__a2bb2o_1 _15949_ (.A1_N(net201),
    .A2_N(net176),
    .B1(_07047_),
    .B2(net155),
    .X(_07050_));
 sky130_fd_sc_hd__o21ai_1 _15950_ (.A1(_06645_),
    .A2(_07049_),
    .B1(_07050_),
    .Y(_07052_));
 sky130_fd_sc_hd__nand2_1 _15951_ (.A(net147),
    .B(_06935_),
    .Y(_07053_));
 sky130_fd_sc_hd__or2_1 _15952_ (.A(_07052_),
    .B(_07053_),
    .X(_07054_));
 sky130_fd_sc_hd__nand2_1 _15953_ (.A(_07052_),
    .B(_07053_),
    .Y(_07055_));
 sky130_fd_sc_hd__and2_2 _15954_ (.A(_07054_),
    .B(_07055_),
    .X(_07056_));
 sky130_fd_sc_hd__nor2_2 _15955_ (.A(net189),
    .B(_06465_),
    .Y(_07057_));
 sky130_fd_sc_hd__nor2_1 _15956_ (.A(_06305_),
    .B(net187),
    .Y(_07058_));
 sky130_fd_sc_hd__o21ba_1 _15957_ (.A1(net189),
    .A2(net134),
    .B1_N(_07058_),
    .X(_07059_));
 sky130_fd_sc_hd__a21o_4 _15958_ (.A1(_06944_),
    .A2(_07057_),
    .B1(_07059_),
    .X(_07060_));
 sky130_fd_sc_hd__nand2_4 _15959_ (.A(net136),
    .B(net184),
    .Y(_07061_));
 sky130_fd_sc_hd__xnor2_4 _15960_ (.A(_07060_),
    .B(_07061_),
    .Y(_07063_));
 sky130_fd_sc_hd__o21a_2 _15961_ (.A1(_06946_),
    .A2(_06947_),
    .B1(_06945_),
    .X(_07064_));
 sky130_fd_sc_hd__nor2_1 _15962_ (.A(_07063_),
    .B(_07064_),
    .Y(_07065_));
 sky130_fd_sc_hd__xor2_4 _15963_ (.A(_07063_),
    .B(_07064_),
    .X(_07066_));
 sky130_fd_sc_hd__xnor2_2 _15964_ (.A(_07056_),
    .B(_07066_),
    .Y(_07067_));
 sky130_fd_sc_hd__a21oi_2 _15965_ (.A1(_06924_),
    .A2(_06926_),
    .B1(_07067_),
    .Y(_07068_));
 sky130_fd_sc_hd__and3_1 _15966_ (.A(_06924_),
    .B(_06926_),
    .C(_07067_),
    .X(_07069_));
 sky130_fd_sc_hd__nor2_1 _15967_ (.A(_07068_),
    .B(_07069_),
    .Y(_07070_));
 sky130_fd_sc_hd__and2_1 _15968_ (.A(_07046_),
    .B(_07070_),
    .X(_07071_));
 sky130_fd_sc_hd__nor2_1 _15969_ (.A(_07046_),
    .B(_07070_),
    .Y(_07072_));
 sky130_fd_sc_hd__or2_2 _15970_ (.A(_07071_),
    .B(_07072_),
    .X(_07074_));
 sky130_fd_sc_hd__nor2_4 _15971_ (.A(_07045_),
    .B(_07074_),
    .Y(_07075_));
 sky130_fd_sc_hd__and2_1 _15972_ (.A(_07045_),
    .B(_07074_),
    .X(_07076_));
 sky130_fd_sc_hd__nor2_4 _15973_ (.A(_07075_),
    .B(_07076_),
    .Y(_07077_));
 sky130_fd_sc_hd__a21oi_4 _15974_ (.A1(_06932_),
    .A2(_06957_),
    .B1(_06930_),
    .Y(_07078_));
 sky130_fd_sc_hd__nand2b_1 _15975_ (.A_N(_07078_),
    .B(_07077_),
    .Y(_07079_));
 sky130_fd_sc_hd__xnor2_4 _15976_ (.A(_07077_),
    .B(_07078_),
    .Y(_07080_));
 sky130_fd_sc_hd__a31o_1 _15977_ (.A1(net147),
    .A2(_06827_),
    .A3(_06940_),
    .B1(_06938_),
    .X(_07081_));
 sky130_fd_sc_hd__o21a_1 _15978_ (.A1(_06954_),
    .A2(_06956_),
    .B1(_07081_),
    .X(_07082_));
 sky130_fd_sc_hd__o21ai_1 _15979_ (.A1(_06954_),
    .A2(_06956_),
    .B1(_07081_),
    .Y(_07083_));
 sky130_fd_sc_hd__nor3_2 _15980_ (.A(_06954_),
    .B(_06956_),
    .C(_07081_),
    .Y(_07085_));
 sky130_fd_sc_hd__nor2_2 _15981_ (.A(_07082_),
    .B(_07085_),
    .Y(_07086_));
 sky130_fd_sc_hd__nand2_4 _15982_ (.A(net142),
    .B(_06827_),
    .Y(_07087_));
 sky130_fd_sc_hd__xnor2_4 _15983_ (.A(_07086_),
    .B(_07087_),
    .Y(_07088_));
 sky130_fd_sc_hd__xnor2_2 _15984_ (.A(_07080_),
    .B(_07088_),
    .Y(_07089_));
 sky130_fd_sc_hd__a21bo_1 _15985_ (.A1(_06960_),
    .A2(_06969_),
    .B1_N(_06959_),
    .X(_07090_));
 sky130_fd_sc_hd__and2b_2 _15986_ (.A_N(_07089_),
    .B(_07090_),
    .X(_07091_));
 sky130_fd_sc_hd__xor2_1 _15987_ (.A(_07089_),
    .B(_07090_),
    .X(_07092_));
 sky130_fd_sc_hd__o21ba_2 _15988_ (.A1(_06965_),
    .A2(_06967_),
    .B1_N(_07092_),
    .X(_07093_));
 sky130_fd_sc_hd__or3b_1 _15989_ (.A(_06965_),
    .B(_06967_),
    .C_N(_07092_),
    .X(_07094_));
 sky130_fd_sc_hd__nand2b_1 _15990_ (.A_N(_07093_),
    .B(_07094_),
    .Y(_07096_));
 sky130_fd_sc_hd__o21ba_2 _15991_ (.A1(_06971_),
    .A2(_06976_),
    .B1_N(_07096_),
    .X(_07097_));
 sky130_fd_sc_hd__or3b_1 _15992_ (.A(_06971_),
    .B(_06976_),
    .C_N(_07096_),
    .X(_07098_));
 sky130_fd_sc_hd__and2b_2 _15993_ (.A_N(_07097_),
    .B(_07098_),
    .X(_07099_));
 sky130_fd_sc_hd__and2_2 _15994_ (.A(_07006_),
    .B(_07098_),
    .X(_07100_));
 sky130_fd_sc_hd__a21oi_2 _15995_ (.A1(_07006_),
    .A2(_07099_),
    .B1(net279),
    .Y(_07101_));
 sky130_fd_sc_hd__o21ai_4 _15996_ (.A1(_07006_),
    .A2(_07099_),
    .B1(_07101_),
    .Y(_07102_));
 sky130_fd_sc_hd__nor2_1 _15997_ (.A(_02260_),
    .B(_02501_),
    .Y(_07103_));
 sky130_fd_sc_hd__or3b_4 _15998_ (.A(net256),
    .B(_07103_),
    .C_N(_02502_),
    .X(_07104_));
 sky130_fd_sc_hd__a21bo_2 _15999_ (.A1(net461),
    .A2(net273),
    .B1_N(net775),
    .X(_07105_));
 sky130_fd_sc_hd__or3b_1 _16000_ (.A(net775),
    .B(net270),
    .C_N(net462),
    .X(_07107_));
 sky130_fd_sc_hd__nand2_1 _16001_ (.A(_07105_),
    .B(_07107_),
    .Y(_07108_));
 sky130_fd_sc_hd__a21boi_2 _16002_ (.A1(_06988_),
    .A2(_06989_),
    .B1_N(_06987_),
    .Y(_07109_));
 sky130_fd_sc_hd__or2_2 _16003_ (.A(_07108_),
    .B(_07109_),
    .X(_07110_));
 sky130_fd_sc_hd__xnor2_1 _16004_ (.A(_07108_),
    .B(_07109_),
    .Y(_07111_));
 sky130_fd_sc_hd__and3_1 _16005_ (.A(_08626_),
    .B(_05780_),
    .C(_05814_),
    .X(_07112_));
 sky130_fd_sc_hd__a21oi_1 _16006_ (.A1(_08626_),
    .A2(_05780_),
    .B1(_05814_),
    .Y(_07113_));
 sky130_fd_sc_hd__or3_1 _16007_ (.A(net252),
    .B(_07112_),
    .C(_07113_),
    .X(_07114_));
 sky130_fd_sc_hd__a221o_1 _16008_ (.A1(_05780_),
    .A2(net239),
    .B1(net234),
    .B2(net774),
    .C1(net243),
    .X(_07115_));
 sky130_fd_sc_hd__o21ba_1 _16009_ (.A1(_08626_),
    .A2(_05945_),
    .B1_N(_07115_),
    .X(_07116_));
 sky130_fd_sc_hd__mux4_2 _16010_ (.A0(_06056_),
    .A1(_06059_),
    .A2(_06061_),
    .A3(_06081_),
    .S0(net297),
    .S1(net302),
    .X(_07118_));
 sky130_fd_sc_hd__or3_1 _16011_ (.A(net569),
    .B(net585),
    .C(_06054_),
    .X(_07119_));
 sky130_fd_sc_hd__mux2_1 _16012_ (.A0(_07118_),
    .A1(_07119_),
    .S(net552),
    .X(_07120_));
 sky130_fd_sc_hd__o22a_1 _16013_ (.A1(net209),
    .A2(_04526_),
    .B1(_05937_),
    .B2(_07120_),
    .X(_07121_));
 sky130_fd_sc_hd__nor2_1 _16014_ (.A(net775),
    .B(_05863_),
    .Y(_07122_));
 sky130_fd_sc_hd__or3_1 _16015_ (.A(net250),
    .B(_05864_),
    .C(_07122_),
    .X(_07123_));
 sky130_fd_sc_hd__o211a_1 _16016_ (.A1(net229),
    .A2(_07111_),
    .B1(_07114_),
    .C1(_07123_),
    .X(_07124_));
 sky130_fd_sc_hd__and3_1 _16017_ (.A(_07116_),
    .B(_07121_),
    .C(_07124_),
    .X(_07125_));
 sky130_fd_sc_hd__a32o_1 _16018_ (.A1(_07102_),
    .A2(_07104_),
    .A3(_07125_),
    .B1(net247),
    .B2(net775),
    .X(_07126_));
 sky130_fd_sc_hd__clkinv_2 _16019_ (.A(_07126_),
    .Y(_08689_));
 sky130_fd_sc_hd__and2_4 _16020_ (.A(net452),
    .B(net226),
    .X(_07128_));
 sky130_fd_sc_hd__nand2_2 _16021_ (.A(net452),
    .B(net227),
    .Y(_07129_));
 sky130_fd_sc_hd__a22o_2 _16022_ (.A1(net140),
    .A2(_06827_),
    .B1(_07128_),
    .B2(_05919_),
    .X(_07130_));
 sky130_fd_sc_hd__nand2_2 _16023_ (.A(net797),
    .B(_07128_),
    .Y(_07131_));
 sky130_fd_sc_hd__o21ai_4 _16024_ (.A1(_06099_),
    .A2(_07131_),
    .B1(_07130_),
    .Y(_07132_));
 sky130_fd_sc_hd__nor2_2 _16025_ (.A(_05987_),
    .B(_07009_),
    .Y(_07133_));
 sky130_fd_sc_hd__xnor2_4 _16026_ (.A(_07132_),
    .B(_07133_),
    .Y(_07134_));
 sky130_fd_sc_hd__nand2_1 _16027_ (.A(_07011_),
    .B(_07134_),
    .Y(_07135_));
 sky130_fd_sc_hd__xnor2_4 _16028_ (.A(_07011_),
    .B(_07134_),
    .Y(_07136_));
 sky130_fd_sc_hd__o21a_1 _16029_ (.A1(net138),
    .A2(_06806_),
    .B1(_07015_),
    .X(_07137_));
 sky130_fd_sc_hd__nor2_1 _16030_ (.A(net138),
    .B(_06907_),
    .Y(_07139_));
 sky130_fd_sc_hd__and3_1 _16031_ (.A(net143),
    .B(_06805_),
    .C(_07139_),
    .X(_07140_));
 sky130_fd_sc_hd__or2_4 _16032_ (.A(_07137_),
    .B(_07140_),
    .X(_07141_));
 sky130_fd_sc_hd__nand2_4 _16033_ (.A(net199),
    .B(net224),
    .Y(_07142_));
 sky130_fd_sc_hd__xnor2_4 _16034_ (.A(_07141_),
    .B(_07142_),
    .Y(_07143_));
 sky130_fd_sc_hd__xor2_4 _16035_ (.A(_07136_),
    .B(_07143_),
    .X(_07144_));
 sky130_fd_sc_hd__xnor2_2 _16036_ (.A(_07021_),
    .B(_07144_),
    .Y(_07145_));
 sky130_fd_sc_hd__o31a_2 _16037_ (.A1(net191),
    .A2(_06448_),
    .A3(_07033_),
    .B1(_07032_),
    .X(_07146_));
 sky130_fd_sc_hd__a31o_4 _16038_ (.A1(_06103_),
    .A2(net224),
    .A3(_07014_),
    .B1(_07016_),
    .X(_07147_));
 sky130_fd_sc_hd__nor2_4 _16039_ (.A(net191),
    .B(net186),
    .Y(_07148_));
 sky130_fd_sc_hd__xnor2_1 _16040_ (.A(_07031_),
    .B(_07148_),
    .Y(_07150_));
 sky130_fd_sc_hd__or3_1 _16041_ (.A(net134),
    .B(_06448_),
    .C(_07150_),
    .X(_07151_));
 sky130_fd_sc_hd__o21ai_1 _16042_ (.A1(net134),
    .A2(_06448_),
    .B1(_07150_),
    .Y(_07152_));
 sky130_fd_sc_hd__and2_2 _16043_ (.A(_07151_),
    .B(_07152_),
    .X(_07153_));
 sky130_fd_sc_hd__xor2_4 _16044_ (.A(_07147_),
    .B(_07153_),
    .X(_07154_));
 sky130_fd_sc_hd__and2b_1 _16045_ (.A_N(_07146_),
    .B(_07154_),
    .X(_07155_));
 sky130_fd_sc_hd__xnor2_2 _16046_ (.A(_07146_),
    .B(_07154_),
    .Y(_07156_));
 sky130_fd_sc_hd__and2b_1 _16047_ (.A_N(_07145_),
    .B(_07156_),
    .X(_07157_));
 sky130_fd_sc_hd__xnor2_2 _16048_ (.A(_07145_),
    .B(_07156_),
    .Y(_07158_));
 sky130_fd_sc_hd__a21oi_2 _16049_ (.A1(_07025_),
    .A2(_07041_),
    .B1(_07024_),
    .Y(_07159_));
 sky130_fd_sc_hd__and2b_1 _16050_ (.A_N(_07159_),
    .B(_07158_),
    .X(_07161_));
 sky130_fd_sc_hd__xnor2_1 _16051_ (.A(_07158_),
    .B(_07159_),
    .Y(_07162_));
 sky130_fd_sc_hd__a21oi_2 _16052_ (.A1(_07056_),
    .A2(_07066_),
    .B1(_07065_),
    .Y(_07163_));
 sky130_fd_sc_hd__and2_4 _16053_ (.A(net762),
    .B(net225),
    .X(_07164_));
 sky130_fd_sc_hd__nand2_4 _16054_ (.A(net765),
    .B(net225),
    .Y(_07165_));
 sky130_fd_sc_hd__nor2_4 _16055_ (.A(net201),
    .B(_07165_),
    .Y(_07166_));
 sky130_fd_sc_hd__and3_1 _16056_ (.A(net155),
    .B(_06732_),
    .C(_07166_),
    .X(_07167_));
 sky130_fd_sc_hd__o22a_1 _16057_ (.A1(net201),
    .A2(_06733_),
    .B1(_07165_),
    .B2(_05901_),
    .X(_07168_));
 sky130_fd_sc_hd__nor2_2 _16058_ (.A(_07167_),
    .B(_07168_),
    .Y(_07169_));
 sky130_fd_sc_hd__nand2_1 _16059_ (.A(net147),
    .B(_07047_),
    .Y(_07170_));
 sky130_fd_sc_hd__xor2_2 _16060_ (.A(_07169_),
    .B(_07170_),
    .X(_07172_));
 sky130_fd_sc_hd__nand2_1 _16061_ (.A(net194),
    .B(net184),
    .Y(_07173_));
 sky130_fd_sc_hd__and3_2 _16062_ (.A(_06372_),
    .B(net184),
    .C(_07058_),
    .X(_07174_));
 sky130_fd_sc_hd__and2b_1 _16063_ (.A_N(_07057_),
    .B(_07173_),
    .X(_07175_));
 sky130_fd_sc_hd__nor2_4 _16064_ (.A(_07174_),
    .B(_07175_),
    .Y(_07176_));
 sky130_fd_sc_hd__nand2_2 _16065_ (.A(net136),
    .B(net178),
    .Y(_07177_));
 sky130_fd_sc_hd__xnor2_4 _16066_ (.A(_07176_),
    .B(_07177_),
    .Y(_07178_));
 sky130_fd_sc_hd__o2bb2ai_4 _16067_ (.A1_N(_06944_),
    .A2_N(_07057_),
    .B1(_07060_),
    .B2(_07061_),
    .Y(_07179_));
 sky130_fd_sc_hd__xor2_2 _16068_ (.A(_07178_),
    .B(_07179_),
    .X(_07180_));
 sky130_fd_sc_hd__nand2b_1 _16069_ (.A_N(_07172_),
    .B(_07180_),
    .Y(_07181_));
 sky130_fd_sc_hd__xnor2_1 _16070_ (.A(_07172_),
    .B(_07180_),
    .Y(_07183_));
 sky130_fd_sc_hd__o21a_2 _16071_ (.A1(_07036_),
    .A2(_07038_),
    .B1(_07183_),
    .X(_07184_));
 sky130_fd_sc_hd__nor3_1 _16072_ (.A(_07036_),
    .B(_07038_),
    .C(_07183_),
    .Y(_07185_));
 sky130_fd_sc_hd__nor2_1 _16073_ (.A(_07184_),
    .B(_07185_),
    .Y(_07186_));
 sky130_fd_sc_hd__and2b_1 _16074_ (.A_N(_07163_),
    .B(_07186_),
    .X(_07187_));
 sky130_fd_sc_hd__xnor2_1 _16075_ (.A(_07163_),
    .B(_07186_),
    .Y(_07188_));
 sky130_fd_sc_hd__and2_1 _16076_ (.A(_07162_),
    .B(_07188_),
    .X(_07189_));
 sky130_fd_sc_hd__nor2_1 _16077_ (.A(_07162_),
    .B(_07188_),
    .Y(_07190_));
 sky130_fd_sc_hd__nor2_2 _16078_ (.A(_07189_),
    .B(_07190_),
    .Y(_07191_));
 sky130_fd_sc_hd__o21ai_4 _16079_ (.A1(_07044_),
    .A2(_07075_),
    .B1(_07191_),
    .Y(_07192_));
 sky130_fd_sc_hd__or3_2 _16080_ (.A(_07044_),
    .B(_07075_),
    .C(_07191_),
    .X(_07194_));
 sky130_fd_sc_hd__nand2_4 _16081_ (.A(_07192_),
    .B(_07194_),
    .Y(_07195_));
 sky130_fd_sc_hd__o21a_1 _16082_ (.A1(_06645_),
    .A2(_07049_),
    .B1(_07054_),
    .X(_07196_));
 sky130_fd_sc_hd__o21ba_1 _16083_ (.A1(_07068_),
    .A2(_07071_),
    .B1_N(_07196_),
    .X(_07197_));
 sky130_fd_sc_hd__or3b_1 _16084_ (.A(_07068_),
    .B(_07071_),
    .C_N(_07196_),
    .X(_07198_));
 sky130_fd_sc_hd__and2b_1 _16085_ (.A_N(_07197_),
    .B(_07198_),
    .X(_07199_));
 sky130_fd_sc_hd__and3_1 _16086_ (.A(net142),
    .B(_06935_),
    .C(_07199_),
    .X(_07200_));
 sky130_fd_sc_hd__a21oi_1 _16087_ (.A1(net142),
    .A2(_06935_),
    .B1(_07199_),
    .Y(_07201_));
 sky130_fd_sc_hd__or2_4 _16088_ (.A(_07200_),
    .B(_07201_),
    .X(_07202_));
 sky130_fd_sc_hd__xnor2_4 _16089_ (.A(_07195_),
    .B(_07202_),
    .Y(_07203_));
 sky130_fd_sc_hd__a21bo_4 _16090_ (.A1(_07080_),
    .A2(_07088_),
    .B1_N(_07079_),
    .X(_07205_));
 sky130_fd_sc_hd__nand2b_1 _16091_ (.A_N(_07203_),
    .B(_07205_),
    .Y(_07206_));
 sky130_fd_sc_hd__xnor2_4 _16092_ (.A(_07203_),
    .B(_07205_),
    .Y(_07207_));
 sky130_fd_sc_hd__o21a_2 _16093_ (.A1(_07085_),
    .A2(_07087_),
    .B1(_07083_),
    .X(_07208_));
 sky130_fd_sc_hd__nand2b_1 _16094_ (.A_N(_07208_),
    .B(_07207_),
    .Y(_07209_));
 sky130_fd_sc_hd__xnor2_4 _16095_ (.A(_07207_),
    .B(_07208_),
    .Y(_07210_));
 sky130_fd_sc_hd__nor3_2 _16096_ (.A(_07091_),
    .B(_07093_),
    .C(_07210_),
    .Y(_07211_));
 sky130_fd_sc_hd__o21ai_4 _16097_ (.A1(_07091_),
    .A2(_07093_),
    .B1(_07210_),
    .Y(_07212_));
 sky130_fd_sc_hd__clkinv_2 _16098_ (.A(_07212_),
    .Y(_07213_));
 sky130_fd_sc_hd__a211o_1 _16099_ (.A1(_07006_),
    .A2(_07098_),
    .B1(_07213_),
    .C1(_07097_),
    .X(_07214_));
 sky130_fd_sc_hd__nor2_1 _16100_ (.A(_07211_),
    .B(_07213_),
    .Y(_07216_));
 sky130_fd_sc_hd__o21bai_4 _16101_ (.A1(_07097_),
    .A2(_07100_),
    .B1_N(_07211_),
    .Y(_07217_));
 sky130_fd_sc_hd__o31a_1 _16102_ (.A1(_07097_),
    .A2(_07100_),
    .A3(_07216_),
    .B1(net281),
    .X(_07218_));
 sky130_fd_sc_hd__o21ai_4 _16103_ (.A1(_07213_),
    .A2(_07217_),
    .B1(_07218_),
    .Y(_07219_));
 sky130_fd_sc_hd__o21ai_4 _16104_ (.A1(_02257_),
    .A2(_02259_),
    .B1(_02502_),
    .Y(_07220_));
 sky130_fd_sc_hd__xor2_4 _16105_ (.A(_02503_),
    .B(_07220_),
    .X(_07221_));
 sky130_fd_sc_hd__nand2_1 _16106_ (.A(net261),
    .B(_07221_),
    .Y(_07222_));
 sky130_fd_sc_hd__a21boi_4 _16107_ (.A1(net453),
    .A2(net273),
    .B1_N(net764),
    .Y(_07223_));
 sky130_fd_sc_hd__and3b_2 _16108_ (.A_N(net764),
    .B(net275),
    .C(net451),
    .X(_07224_));
 sky130_fd_sc_hd__a211oi_4 _16109_ (.A1(_07105_),
    .A2(_07110_),
    .B1(_07223_),
    .C1(_07224_),
    .Y(_07225_));
 sky130_fd_sc_hd__o211a_1 _16110_ (.A1(_07223_),
    .A2(_07224_),
    .B1(_07105_),
    .C1(_07110_),
    .X(_07227_));
 sky130_fd_sc_hd__or3_1 _16111_ (.A(net228),
    .B(_07225_),
    .C(_07227_),
    .X(_07228_));
 sky130_fd_sc_hd__and3_1 _16112_ (.A(_05001_),
    .B(_05778_),
    .C(_05815_),
    .X(_07229_));
 sky130_fd_sc_hd__a21oi_1 _16113_ (.A1(_05001_),
    .A2(_05778_),
    .B1(_05815_),
    .Y(_07230_));
 sky130_fd_sc_hd__nor2_1 _16114_ (.A(net764),
    .B(_05864_),
    .Y(_07231_));
 sky130_fd_sc_hd__or3_1 _16115_ (.A(net251),
    .B(_05865_),
    .C(_07231_),
    .X(_07232_));
 sky130_fd_sc_hd__mux4_2 _16116_ (.A0(_06124_),
    .A1(_06128_),
    .A2(_06130_),
    .A3(_06153_),
    .S0(net299),
    .S1(net303),
    .X(_07233_));
 sky130_fd_sc_hd__o31a_1 _16117_ (.A1(net577),
    .A2(net592),
    .A3(_06122_),
    .B1(net559),
    .X(_07234_));
 sky130_fd_sc_hd__a211o_1 _16118_ (.A1(_03203_),
    .A2(_07233_),
    .B1(_07234_),
    .C1(net241),
    .X(_07235_));
 sky130_fd_sc_hd__a221o_1 _16119_ (.A1(_05778_),
    .A2(net239),
    .B1(net233),
    .B2(net764),
    .C1(net244),
    .X(_07236_));
 sky130_fd_sc_hd__a31o_1 _16120_ (.A1(net451),
    .A2(net764),
    .A3(net236),
    .B1(_07236_),
    .X(_07238_));
 sky130_fd_sc_hd__a21oi_1 _16121_ (.A1(_02643_),
    .A2(_04754_),
    .B1(_07238_),
    .Y(_07239_));
 sky130_fd_sc_hd__and3_1 _16122_ (.A(_07232_),
    .B(_07235_),
    .C(_07239_),
    .X(_07240_));
 sky130_fd_sc_hd__o311a_1 _16123_ (.A1(net253),
    .A2(_07229_),
    .A3(_07230_),
    .B1(_07240_),
    .C1(_07228_),
    .X(_07241_));
 sky130_fd_sc_hd__a32o_1 _16124_ (.A1(_07219_),
    .A2(_07222_),
    .A3(_07241_),
    .B1(net247),
    .B2(net763),
    .X(_07242_));
 sky130_fd_sc_hd__clkinv_2 _16125_ (.A(_07242_),
    .Y(_08690_));
 sky130_fd_sc_hd__o22a_1 _16126_ (.A1(net139),
    .A2(_06936_),
    .B1(_07129_),
    .B2(_05987_),
    .X(_07243_));
 sky130_fd_sc_hd__and3_1 _16127_ (.A(net148),
    .B(net140),
    .C(_07128_),
    .X(_07244_));
 sky130_fd_sc_hd__a21o_2 _16128_ (.A1(net784),
    .A2(_07244_),
    .B1(_07243_),
    .X(_07245_));
 sky130_fd_sc_hd__nand2_2 _16129_ (.A(net143),
    .B(_07008_),
    .Y(_07246_));
 sky130_fd_sc_hd__xor2_4 _16130_ (.A(_07245_),
    .B(_07246_),
    .X(_07248_));
 sky130_fd_sc_hd__a2bb2o_2 _16131_ (.A1_N(_06099_),
    .A2_N(_07131_),
    .B1(_07133_),
    .B2(_07130_),
    .X(_07249_));
 sky130_fd_sc_hd__and2_1 _16132_ (.A(_07248_),
    .B(_07249_),
    .X(_07250_));
 sky130_fd_sc_hd__xnor2_2 _16133_ (.A(_07248_),
    .B(_07249_),
    .Y(_07251_));
 sky130_fd_sc_hd__nand2_1 _16134_ (.A(net480),
    .B(net198),
    .Y(_07252_));
 sky130_fd_sc_hd__o21a_1 _16135_ (.A1(net138),
    .A2(_06907_),
    .B1(_07252_),
    .X(_07253_));
 sky130_fd_sc_hd__and3_1 _16136_ (.A(net480),
    .B(net199),
    .C(_07139_),
    .X(_07254_));
 sky130_fd_sc_hd__or2_2 _16137_ (.A(_07253_),
    .B(_07254_),
    .X(_07255_));
 sky130_fd_sc_hd__nor2_2 _16138_ (.A(_06247_),
    .B(_06712_),
    .Y(_07256_));
 sky130_fd_sc_hd__and2b_1 _16139_ (.A_N(_07255_),
    .B(_07256_),
    .X(_07257_));
 sky130_fd_sc_hd__xor2_2 _16140_ (.A(_07255_),
    .B(_07256_),
    .X(_07259_));
 sky130_fd_sc_hd__nor2_2 _16141_ (.A(_07251_),
    .B(_07259_),
    .Y(_07260_));
 sky130_fd_sc_hd__and2_1 _16142_ (.A(_07251_),
    .B(_07259_),
    .X(_07261_));
 sky130_fd_sc_hd__nor2_4 _16143_ (.A(_07260_),
    .B(_07261_),
    .Y(_07262_));
 sky130_fd_sc_hd__o21a_2 _16144_ (.A1(_07136_),
    .A2(_07143_),
    .B1(_07135_),
    .X(_07263_));
 sky130_fd_sc_hd__nand2b_1 _16145_ (.A_N(_07263_),
    .B(_07262_),
    .Y(_07264_));
 sky130_fd_sc_hd__xnor2_4 _16146_ (.A(_07262_),
    .B(_07263_),
    .Y(_07265_));
 sky130_fd_sc_hd__a21bo_4 _16147_ (.A1(_07031_),
    .A2(_07148_),
    .B1_N(_07151_),
    .X(_07266_));
 sky130_fd_sc_hd__o21ba_4 _16148_ (.A1(_07137_),
    .A2(_07142_),
    .B1_N(_07140_),
    .X(_07267_));
 sky130_fd_sc_hd__o22a_2 _16149_ (.A1(net134),
    .A2(net186),
    .B1(net180),
    .B2(net191),
    .X(_07268_));
 sky130_fd_sc_hd__nor2_4 _16150_ (.A(net134),
    .B(net180),
    .Y(_07270_));
 sky130_fd_sc_hd__a21oi_4 _16151_ (.A1(_07148_),
    .A2(_07270_),
    .B1(_07268_),
    .Y(_07271_));
 sky130_fd_sc_hd__nand2_4 _16152_ (.A(_06447_),
    .B(net188),
    .Y(_07272_));
 sky130_fd_sc_hd__xor2_4 _16153_ (.A(_07271_),
    .B(_07272_),
    .X(_07273_));
 sky130_fd_sc_hd__nor2_1 _16154_ (.A(_07267_),
    .B(_07273_),
    .Y(_07274_));
 sky130_fd_sc_hd__xnor2_4 _16155_ (.A(_07267_),
    .B(_07273_),
    .Y(_07275_));
 sky130_fd_sc_hd__and2b_1 _16156_ (.A_N(_07275_),
    .B(_07266_),
    .X(_07276_));
 sky130_fd_sc_hd__xnor2_4 _16157_ (.A(_07266_),
    .B(_07275_),
    .Y(_07277_));
 sky130_fd_sc_hd__xnor2_4 _16158_ (.A(_07265_),
    .B(_07277_),
    .Y(_07278_));
 sky130_fd_sc_hd__a21oi_4 _16159_ (.A1(_07021_),
    .A2(_07144_),
    .B1(_07157_),
    .Y(_07279_));
 sky130_fd_sc_hd__or2_1 _16160_ (.A(_07278_),
    .B(_07279_),
    .X(_07281_));
 sky130_fd_sc_hd__xnor2_4 _16161_ (.A(_07278_),
    .B(_07279_),
    .Y(_07282_));
 sky130_fd_sc_hd__a21bo_1 _16162_ (.A1(_07178_),
    .A2(_07179_),
    .B1_N(_07181_),
    .X(_07283_));
 sky130_fd_sc_hd__a21oi_2 _16163_ (.A1(_07147_),
    .A2(_07153_),
    .B1(_07155_),
    .Y(_07284_));
 sky130_fd_sc_hd__nand2_1 _16164_ (.A(net147),
    .B(_07164_),
    .Y(_07285_));
 sky130_fd_sc_hd__and3_2 _16165_ (.A(net147),
    .B(_06827_),
    .C(_07166_),
    .X(_07286_));
 sky130_fd_sc_hd__a21oi_4 _16166_ (.A1(_06829_),
    .A2(_07285_),
    .B1(_07286_),
    .Y(_07287_));
 sky130_fd_sc_hd__nor2_1 _16167_ (.A(net189),
    .B(net176),
    .Y(_07288_));
 sky130_fd_sc_hd__or3_4 _16168_ (.A(net189),
    .B(net176),
    .C(_07173_),
    .X(_07289_));
 sky130_fd_sc_hd__a22o_1 _16169_ (.A1(_06372_),
    .A2(net184),
    .B1(net178),
    .B2(net194),
    .X(_07290_));
 sky130_fd_sc_hd__nand2_4 _16170_ (.A(_07289_),
    .B(_07290_),
    .Y(_07292_));
 sky130_fd_sc_hd__nand2_4 _16171_ (.A(net136),
    .B(_06732_),
    .Y(_07293_));
 sky130_fd_sc_hd__xor2_4 _16172_ (.A(_07292_),
    .B(_07293_),
    .X(_07294_));
 sky130_fd_sc_hd__a31o_4 _16173_ (.A1(net137),
    .A2(net178),
    .A3(_07176_),
    .B1(_07174_),
    .X(_07295_));
 sky130_fd_sc_hd__xor2_4 _16174_ (.A(_07294_),
    .B(_07295_),
    .X(_07296_));
 sky130_fd_sc_hd__xor2_2 _16175_ (.A(_07287_),
    .B(_07296_),
    .X(_07297_));
 sky130_fd_sc_hd__and2b_1 _16176_ (.A_N(_07284_),
    .B(_07297_),
    .X(_07298_));
 sky130_fd_sc_hd__xnor2_1 _16177_ (.A(_07284_),
    .B(_07297_),
    .Y(_07299_));
 sky130_fd_sc_hd__and2_2 _16178_ (.A(_07283_),
    .B(_07299_),
    .X(_07300_));
 sky130_fd_sc_hd__nor2_1 _16179_ (.A(_07283_),
    .B(_07299_),
    .Y(_07301_));
 sky130_fd_sc_hd__nor2_1 _16180_ (.A(_07300_),
    .B(_07301_),
    .Y(_07303_));
 sky130_fd_sc_hd__xnor2_2 _16181_ (.A(_07282_),
    .B(_07303_),
    .Y(_07304_));
 sky130_fd_sc_hd__o21a_1 _16182_ (.A1(_07161_),
    .A2(_07189_),
    .B1(_07304_),
    .X(_07305_));
 sky130_fd_sc_hd__nor3_1 _16183_ (.A(_07161_),
    .B(_07189_),
    .C(_07304_),
    .Y(_07306_));
 sky130_fd_sc_hd__nor2_2 _16184_ (.A(_07305_),
    .B(_07306_),
    .Y(_07307_));
 sky130_fd_sc_hd__a31o_2 _16185_ (.A1(net147),
    .A2(_07047_),
    .A3(_07169_),
    .B1(_07167_),
    .X(_07308_));
 sky130_fd_sc_hd__o21a_1 _16186_ (.A1(_07184_),
    .A2(_07187_),
    .B1(_07308_),
    .X(_07309_));
 sky130_fd_sc_hd__o21ai_1 _16187_ (.A1(_07184_),
    .A2(_07187_),
    .B1(_07308_),
    .Y(_07310_));
 sky130_fd_sc_hd__nor3_2 _16188_ (.A(_07184_),
    .B(_07187_),
    .C(_07308_),
    .Y(_07311_));
 sky130_fd_sc_hd__nor2_2 _16189_ (.A(_07309_),
    .B(_07311_),
    .Y(_07312_));
 sky130_fd_sc_hd__nand2_4 _16190_ (.A(net142),
    .B(_07047_),
    .Y(_07314_));
 sky130_fd_sc_hd__xnor2_4 _16191_ (.A(_07312_),
    .B(_07314_),
    .Y(_07315_));
 sky130_fd_sc_hd__xnor2_2 _16192_ (.A(_07307_),
    .B(_07315_),
    .Y(_07316_));
 sky130_fd_sc_hd__o21a_1 _16193_ (.A1(_07195_),
    .A2(_07202_),
    .B1(_07192_),
    .X(_07317_));
 sky130_fd_sc_hd__nor2_1 _16194_ (.A(_07316_),
    .B(_07317_),
    .Y(_07318_));
 sky130_fd_sc_hd__xnor2_1 _16195_ (.A(_07316_),
    .B(_07317_),
    .Y(_07319_));
 sky130_fd_sc_hd__o21ba_1 _16196_ (.A1(_07197_),
    .A2(_07200_),
    .B1_N(_07319_),
    .X(_07320_));
 sky130_fd_sc_hd__or3b_1 _16197_ (.A(_07197_),
    .B(_07200_),
    .C_N(_07319_),
    .X(_07321_));
 sky130_fd_sc_hd__nand2b_1 _16198_ (.A_N(_07320_),
    .B(_07321_),
    .Y(_07322_));
 sky130_fd_sc_hd__a21oi_2 _16199_ (.A1(_07206_),
    .A2(_07209_),
    .B1(_07322_),
    .Y(_07323_));
 sky130_fd_sc_hd__and3_1 _16200_ (.A(_07206_),
    .B(_07209_),
    .C(_07322_),
    .X(_07325_));
 sky130_fd_sc_hd__or2_4 _16201_ (.A(_07323_),
    .B(_07325_),
    .X(_07326_));
 sky130_fd_sc_hd__a21oi_4 _16202_ (.A1(_07212_),
    .A2(_07217_),
    .B1(_07326_),
    .Y(_07327_));
 sky130_fd_sc_hd__or3b_4 _16203_ (.A(_07211_),
    .B(_07326_),
    .C_N(_07214_),
    .X(_07328_));
 sky130_fd_sc_hd__a31o_1 _16204_ (.A1(_07212_),
    .A2(_07217_),
    .A3(_07326_),
    .B1(net279),
    .X(_07329_));
 sky130_fd_sc_hd__or2_4 _16205_ (.A(_07327_),
    .B(_07329_),
    .X(_07330_));
 sky130_fd_sc_hd__nor2_1 _16206_ (.A(_02505_),
    .B(_02508_),
    .Y(_07331_));
 sky130_fd_sc_hd__or3_4 _16207_ (.A(_02509_),
    .B(net256),
    .C(_07331_),
    .X(_07332_));
 sky130_fd_sc_hd__a21boi_4 _16208_ (.A1(net444),
    .A2(net273),
    .B1_N(net753),
    .Y(_07333_));
 sky130_fd_sc_hd__and3b_1 _16209_ (.A_N(net753),
    .B(net273),
    .C(net444),
    .X(_07334_));
 sky130_fd_sc_hd__nor2_1 _16210_ (.A(_07333_),
    .B(_07334_),
    .Y(_07336_));
 sky130_fd_sc_hd__o21ba_1 _16211_ (.A1(_07223_),
    .A2(_07225_),
    .B1_N(_07334_),
    .X(_07337_));
 sky130_fd_sc_hd__o21ai_1 _16212_ (.A1(_07223_),
    .A2(_07225_),
    .B1(_07336_),
    .Y(_07338_));
 sky130_fd_sc_hd__o31a_1 _16213_ (.A1(_07223_),
    .A2(_07225_),
    .A3(_07336_),
    .B1(_05951_),
    .X(_07339_));
 sky130_fd_sc_hd__a21oi_1 _16214_ (.A1(_03648_),
    .A2(_05777_),
    .B1(_05816_),
    .Y(_07340_));
 sky130_fd_sc_hd__a311o_1 _16215_ (.A1(_03648_),
    .A2(_05777_),
    .A3(_05816_),
    .B1(net252),
    .C1(_07340_),
    .X(_07341_));
 sky130_fd_sc_hd__a21oi_1 _16216_ (.A1(net753),
    .A2(_05865_),
    .B1(net251),
    .Y(_07342_));
 sky130_fd_sc_hd__o21a_1 _16217_ (.A1(net753),
    .A2(_05865_),
    .B1(_07342_),
    .X(_07343_));
 sky130_fd_sc_hd__a221o_1 _16218_ (.A1(_05777_),
    .A2(net238),
    .B1(net233),
    .B2(net754),
    .C1(net244),
    .X(_07344_));
 sky130_fd_sc_hd__o22ai_2 _16219_ (.A1(net210),
    .A2(_04760_),
    .B1(net203),
    .B2(_05978_),
    .Y(_07345_));
 sky130_fd_sc_hd__a211o_1 _16220_ (.A1(_03637_),
    .A2(net236),
    .B1(_07344_),
    .C1(_07345_),
    .X(_07347_));
 sky130_fd_sc_hd__or3b_2 _16221_ (.A(_07347_),
    .B(_07343_),
    .C_N(_07341_),
    .X(_07348_));
 sky130_fd_sc_hd__a21oi_1 _16222_ (.A1(_07338_),
    .A2(_07339_),
    .B1(_07348_),
    .Y(_07349_));
 sky130_fd_sc_hd__a32o_1 _16223_ (.A1(_07330_),
    .A2(_07332_),
    .A3(_07349_),
    .B1(net247),
    .B2(net753),
    .X(_07350_));
 sky130_fd_sc_hd__clkinv_2 _16224_ (.A(_07350_),
    .Y(_08691_));
 sky130_fd_sc_hd__o22a_1 _16225_ (.A1(net139),
    .A2(_07048_),
    .B1(_07129_),
    .B2(_06042_),
    .X(_07351_));
 sky130_fd_sc_hd__and4_2 _16226_ (.A(net774),
    .B(net143),
    .C(net140),
    .D(_07128_),
    .X(_07352_));
 sky130_fd_sc_hd__nor2_4 _16227_ (.A(_07351_),
    .B(_07352_),
    .Y(_07353_));
 sky130_fd_sc_hd__nor2_4 _16228_ (.A(_06104_),
    .B(_07009_),
    .Y(_07354_));
 sky130_fd_sc_hd__xor2_4 _16229_ (.A(_07353_),
    .B(_07354_),
    .X(_07355_));
 sky130_fd_sc_hd__a2bb2o_2 _16230_ (.A1_N(_07243_),
    .A2_N(_07246_),
    .B1(_07244_),
    .B2(net784),
    .X(_07357_));
 sky130_fd_sc_hd__nand2_1 _16231_ (.A(_07355_),
    .B(_07357_),
    .Y(_07358_));
 sky130_fd_sc_hd__xor2_2 _16232_ (.A(_07355_),
    .B(_07357_),
    .X(_07359_));
 sky130_fd_sc_hd__a22o_1 _16233_ (.A1(net471),
    .A2(net198),
    .B1(net197),
    .B2(_06805_),
    .X(_07360_));
 sky130_fd_sc_hd__or3_1 _16234_ (.A(net196),
    .B(_06907_),
    .C(_07252_),
    .X(_07361_));
 sky130_fd_sc_hd__and2_2 _16235_ (.A(_07360_),
    .B(_07361_),
    .X(_07362_));
 sky130_fd_sc_hd__nor2_2 _16236_ (.A(net191),
    .B(_06712_),
    .Y(_07363_));
 sky130_fd_sc_hd__nand2_1 _16237_ (.A(_07362_),
    .B(_07363_),
    .Y(_07364_));
 sky130_fd_sc_hd__xor2_2 _16238_ (.A(_07362_),
    .B(_07363_),
    .X(_07365_));
 sky130_fd_sc_hd__xnor2_1 _16239_ (.A(_07359_),
    .B(_07365_),
    .Y(_07366_));
 sky130_fd_sc_hd__o21ba_1 _16240_ (.A1(_07250_),
    .A2(_07260_),
    .B1_N(_07366_),
    .X(_07368_));
 sky130_fd_sc_hd__or3b_4 _16241_ (.A(_07250_),
    .B(_07260_),
    .C_N(_07366_),
    .X(_07369_));
 sky130_fd_sc_hd__nand2b_4 _16242_ (.A_N(_07368_),
    .B(_07369_),
    .Y(_07370_));
 sky130_fd_sc_hd__a2bb2o_4 _16243_ (.A1_N(_07268_),
    .A2_N(_07272_),
    .B1(_07270_),
    .B2(_07148_),
    .X(_07371_));
 sky130_fd_sc_hd__nor2_1 _16244_ (.A(_06465_),
    .B(net185),
    .Y(_07372_));
 sky130_fd_sc_hd__xor2_1 _16245_ (.A(_07270_),
    .B(_07372_),
    .X(_07373_));
 sky130_fd_sc_hd__and3_1 _16246_ (.A(net131),
    .B(_06552_),
    .C(_07373_),
    .X(_07374_));
 sky130_fd_sc_hd__a21oi_1 _16247_ (.A1(net131),
    .A2(_06552_),
    .B1(_07373_),
    .Y(_07375_));
 sky130_fd_sc_hd__nor2_1 _16248_ (.A(_07374_),
    .B(_07375_),
    .Y(_07376_));
 sky130_fd_sc_hd__o21a_2 _16249_ (.A1(_07254_),
    .A2(_07257_),
    .B1(_07376_),
    .X(_07377_));
 sky130_fd_sc_hd__nor3_2 _16250_ (.A(_07254_),
    .B(_07257_),
    .C(_07376_),
    .Y(_07379_));
 sky130_fd_sc_hd__nor2_4 _16251_ (.A(_07377_),
    .B(_07379_),
    .Y(_07380_));
 sky130_fd_sc_hd__xnor2_4 _16252_ (.A(_07371_),
    .B(_07380_),
    .Y(_07381_));
 sky130_fd_sc_hd__nor2_1 _16253_ (.A(_07370_),
    .B(_07381_),
    .Y(_07382_));
 sky130_fd_sc_hd__xor2_4 _16254_ (.A(_07370_),
    .B(_07381_),
    .X(_07383_));
 sky130_fd_sc_hd__a21bo_1 _16255_ (.A1(_07265_),
    .A2(_07277_),
    .B1_N(_07264_),
    .X(_07384_));
 sky130_fd_sc_hd__and2_1 _16256_ (.A(_07383_),
    .B(_07384_),
    .X(_07385_));
 sky130_fd_sc_hd__xor2_2 _16257_ (.A(_07383_),
    .B(_07384_),
    .X(_07386_));
 sky130_fd_sc_hd__a22oi_4 _16258_ (.A1(_07294_),
    .A2(_07295_),
    .B1(_07296_),
    .B2(_07287_),
    .Y(_07387_));
 sky130_fd_sc_hd__and3_1 _16259_ (.A(net194),
    .B(net174),
    .C(_07288_),
    .X(_07388_));
 sky130_fd_sc_hd__a21oi_1 _16260_ (.A1(net194),
    .A2(net174),
    .B1(_07288_),
    .Y(_07390_));
 sky130_fd_sc_hd__or2_1 _16261_ (.A(_07388_),
    .B(_07390_),
    .X(_07391_));
 sky130_fd_sc_hd__nor3_2 _16262_ (.A(_06236_),
    .B(_06828_),
    .C(_07391_),
    .Y(_07392_));
 sky130_fd_sc_hd__o21a_1 _16263_ (.A1(_06236_),
    .A2(_06828_),
    .B1(_07391_),
    .X(_07393_));
 sky130_fd_sc_hd__nor2_2 _16264_ (.A(_07392_),
    .B(_07393_),
    .Y(_07394_));
 sky130_fd_sc_hd__o21ai_4 _16265_ (.A1(_07292_),
    .A2(_07293_),
    .B1(_07289_),
    .Y(_07395_));
 sky130_fd_sc_hd__xor2_2 _16266_ (.A(_07394_),
    .B(_07395_),
    .X(_07396_));
 sky130_fd_sc_hd__nand2b_1 _16267_ (.A_N(_06937_),
    .B(_07396_),
    .Y(_07397_));
 sky130_fd_sc_hd__xnor2_1 _16268_ (.A(_06937_),
    .B(_07396_),
    .Y(_07398_));
 sky130_fd_sc_hd__o21a_1 _16269_ (.A1(_07274_),
    .A2(_07276_),
    .B1(_07398_),
    .X(_07399_));
 sky130_fd_sc_hd__nor3_1 _16270_ (.A(_07274_),
    .B(_07276_),
    .C(_07398_),
    .Y(_07401_));
 sky130_fd_sc_hd__nor2_1 _16271_ (.A(_07399_),
    .B(_07401_),
    .Y(_07402_));
 sky130_fd_sc_hd__xnor2_2 _16272_ (.A(_07387_),
    .B(_07402_),
    .Y(_07403_));
 sky130_fd_sc_hd__xnor2_1 _16273_ (.A(_07386_),
    .B(_07403_),
    .Y(_07404_));
 sky130_fd_sc_hd__o31a_1 _16274_ (.A1(_07282_),
    .A2(_07300_),
    .A3(_07301_),
    .B1(_07281_),
    .X(_07405_));
 sky130_fd_sc_hd__or2_2 _16275_ (.A(_07404_),
    .B(_07405_),
    .X(_07406_));
 sky130_fd_sc_hd__nand2_1 _16276_ (.A(_07404_),
    .B(_07405_),
    .Y(_07407_));
 sky130_fd_sc_hd__nand2_4 _16277_ (.A(_07406_),
    .B(_07407_),
    .Y(_07408_));
 sky130_fd_sc_hd__o21a_1 _16278_ (.A1(_07298_),
    .A2(_07300_),
    .B1(_07286_),
    .X(_07409_));
 sky130_fd_sc_hd__nor3_2 _16279_ (.A(_07286_),
    .B(_07298_),
    .C(_07300_),
    .Y(_07410_));
 sky130_fd_sc_hd__nor2_4 _16280_ (.A(_07409_),
    .B(_07410_),
    .Y(_07412_));
 sky130_fd_sc_hd__nand2_4 _16281_ (.A(net142),
    .B(_07164_),
    .Y(_07413_));
 sky130_fd_sc_hd__xor2_4 _16282_ (.A(_07412_),
    .B(_07413_),
    .X(_07414_));
 sky130_fd_sc_hd__xor2_4 _16283_ (.A(_07408_),
    .B(_07414_),
    .X(_07415_));
 sky130_fd_sc_hd__a21o_1 _16284_ (.A1(_07307_),
    .A2(_07315_),
    .B1(_07305_),
    .X(_07416_));
 sky130_fd_sc_hd__xor2_2 _16285_ (.A(_07415_),
    .B(_07416_),
    .X(_07417_));
 sky130_fd_sc_hd__o21a_1 _16286_ (.A1(_07311_),
    .A2(_07314_),
    .B1(_07310_),
    .X(_07418_));
 sky130_fd_sc_hd__nand2b_1 _16287_ (.A_N(_07418_),
    .B(_07417_),
    .Y(_07419_));
 sky130_fd_sc_hd__xnor2_1 _16288_ (.A(_07417_),
    .B(_07418_),
    .Y(_07420_));
 sky130_fd_sc_hd__o21a_1 _16289_ (.A1(_07318_),
    .A2(_07320_),
    .B1(_07420_),
    .X(_07421_));
 sky130_fd_sc_hd__or3_4 _16290_ (.A(_07318_),
    .B(_07320_),
    .C(_07420_),
    .X(_07423_));
 sky130_fd_sc_hd__nand2b_4 _16291_ (.A_N(_07421_),
    .B(_07423_),
    .Y(_07424_));
 sky130_fd_sc_hd__nor2_2 _16292_ (.A(_07323_),
    .B(_07327_),
    .Y(_07425_));
 sky130_fd_sc_hd__xnor2_4 _16293_ (.A(_07424_),
    .B(_07425_),
    .Y(_07426_));
 sky130_fd_sc_hd__nor2_2 _16294_ (.A(_02507_),
    .B(_02509_),
    .Y(_07427_));
 sky130_fd_sc_hd__xnor2_4 _16295_ (.A(_02097_),
    .B(_07427_),
    .Y(_07428_));
 sky130_fd_sc_hd__nand2_2 _16296_ (.A(net261),
    .B(_07428_),
    .Y(_07429_));
 sky130_fd_sc_hd__a21bo_1 _16297_ (.A1(net434),
    .A2(net274),
    .B1_N(net744),
    .X(_07430_));
 sky130_fd_sc_hd__or3b_2 _16298_ (.A(net744),
    .B(net271),
    .C_N(net435),
    .X(_07431_));
 sky130_fd_sc_hd__nand2_1 _16299_ (.A(_07430_),
    .B(_07431_),
    .Y(_07432_));
 sky130_fd_sc_hd__nor2_1 _16300_ (.A(_07333_),
    .B(_07337_),
    .Y(_07434_));
 sky130_fd_sc_hd__xnor2_1 _16301_ (.A(_07432_),
    .B(_07434_),
    .Y(_07435_));
 sky130_fd_sc_hd__and3_1 _16302_ (.A(_03659_),
    .B(_05776_),
    .C(_05817_),
    .X(_07436_));
 sky130_fd_sc_hd__a21oi_1 _16303_ (.A1(_03659_),
    .A2(_05776_),
    .B1(_05817_),
    .Y(_07437_));
 sky130_fd_sc_hd__or3_1 _16304_ (.A(net252),
    .B(_07436_),
    .C(_07437_),
    .X(_07438_));
 sky130_fd_sc_hd__a21oi_1 _16305_ (.A1(net753),
    .A2(_05865_),
    .B1(net744),
    .Y(_07439_));
 sky130_fd_sc_hd__or3_1 _16306_ (.A(net251),
    .B(_05866_),
    .C(_07439_),
    .X(_07440_));
 sky130_fd_sc_hd__a221o_1 _16307_ (.A1(_05776_),
    .A2(net238),
    .B1(net232),
    .B2(net744),
    .C1(net245),
    .X(_07441_));
 sky130_fd_sc_hd__o21ba_1 _16308_ (.A1(_03659_),
    .A2(net235),
    .B1_N(_07441_),
    .X(_07442_));
 sky130_fd_sc_hd__o22a_1 _16309_ (.A1(net210),
    .A2(_04874_),
    .B1(net202),
    .B2(_06009_),
    .X(_07443_));
 sky130_fd_sc_hd__and4_1 _16310_ (.A(_07438_),
    .B(_07440_),
    .C(_07442_),
    .D(_07443_),
    .X(_07445_));
 sky130_fd_sc_hd__o221a_1 _16311_ (.A1(net278),
    .A2(_07426_),
    .B1(_07435_),
    .B2(net229),
    .C1(_07445_),
    .X(_07446_));
 sky130_fd_sc_hd__a22o_1 _16312_ (.A1(net744),
    .A2(net248),
    .B1(_07429_),
    .B2(_07446_),
    .X(_07447_));
 sky130_fd_sc_hd__inv_2 _16313_ (.A(_07447_),
    .Y(_08692_));
 sky130_fd_sc_hd__a22o_1 _16314_ (.A1(_06103_),
    .A2(_07128_),
    .B1(_07164_),
    .B2(net140),
    .X(_07448_));
 sky130_fd_sc_hd__or4_4 _16315_ (.A(_05001_),
    .B(_06098_),
    .C(net138),
    .D(net267),
    .X(_07449_));
 sky130_fd_sc_hd__nand2_4 _16316_ (.A(_07448_),
    .B(_07449_),
    .Y(_07450_));
 sky130_fd_sc_hd__nand2_4 _16317_ (.A(net461),
    .B(net198),
    .Y(_07451_));
 sky130_fd_sc_hd__xnor2_2 _16318_ (.A(_07450_),
    .B(_07451_),
    .Y(_07452_));
 sky130_fd_sc_hd__a21o_1 _16319_ (.A1(_07353_),
    .A2(_07354_),
    .B1(_07352_),
    .X(_07453_));
 sky130_fd_sc_hd__and2b_1 _16320_ (.A_N(_07452_),
    .B(_07453_),
    .X(_07455_));
 sky130_fd_sc_hd__xor2_1 _16321_ (.A(_07452_),
    .B(_07453_),
    .X(_07456_));
 sky130_fd_sc_hd__a22o_1 _16322_ (.A1(_06313_),
    .A2(net172),
    .B1(_06906_),
    .B2(net197),
    .X(_07457_));
 sky130_fd_sc_hd__or4_1 _16323_ (.A(net196),
    .B(net191),
    .C(net171),
    .D(net169),
    .X(_07458_));
 sky130_fd_sc_hd__nand2_1 _16324_ (.A(_07457_),
    .B(_07458_),
    .Y(_07459_));
 sky130_fd_sc_hd__nor2_1 _16325_ (.A(net133),
    .B(_06712_),
    .Y(_07460_));
 sky130_fd_sc_hd__xor2_1 _16326_ (.A(_07459_),
    .B(_07460_),
    .X(_07461_));
 sky130_fd_sc_hd__and2_1 _16327_ (.A(_07456_),
    .B(_07461_),
    .X(_07462_));
 sky130_fd_sc_hd__nor2_1 _16328_ (.A(_07456_),
    .B(_07461_),
    .Y(_07463_));
 sky130_fd_sc_hd__nor2_1 _16329_ (.A(_07462_),
    .B(_07463_),
    .Y(_07464_));
 sky130_fd_sc_hd__a21bo_1 _16330_ (.A1(_07359_),
    .A2(_07365_),
    .B1_N(_07358_),
    .X(_07466_));
 sky130_fd_sc_hd__xor2_1 _16331_ (.A(_07464_),
    .B(_07466_),
    .X(_07467_));
 sky130_fd_sc_hd__a21oi_2 _16332_ (.A1(_07270_),
    .A2(_07372_),
    .B1(_07374_),
    .Y(_07468_));
 sky130_fd_sc_hd__o22a_2 _16333_ (.A1(net185),
    .A2(net183),
    .B1(net179),
    .B2(net187),
    .X(_07469_));
 sky130_fd_sc_hd__or4_4 _16334_ (.A(net187),
    .B(net185),
    .C(net183),
    .D(net179),
    .X(_07470_));
 sky130_fd_sc_hd__nand2b_1 _16335_ (.A_N(_07469_),
    .B(_07470_),
    .Y(_07471_));
 sky130_fd_sc_hd__nand2_2 _16336_ (.A(net132),
    .B(net177),
    .Y(_07472_));
 sky130_fd_sc_hd__xnor2_1 _16337_ (.A(_07471_),
    .B(_07472_),
    .Y(_07473_));
 sky130_fd_sc_hd__a21oi_1 _16338_ (.A1(_07361_),
    .A2(_07364_),
    .B1(_07473_),
    .Y(_07474_));
 sky130_fd_sc_hd__and3_1 _16339_ (.A(_07361_),
    .B(_07364_),
    .C(_07473_),
    .X(_07475_));
 sky130_fd_sc_hd__nor2_1 _16340_ (.A(_07474_),
    .B(_07475_),
    .Y(_07477_));
 sky130_fd_sc_hd__and2b_1 _16341_ (.A_N(_07468_),
    .B(_07477_),
    .X(_07478_));
 sky130_fd_sc_hd__xnor2_1 _16342_ (.A(_07468_),
    .B(_07477_),
    .Y(_07479_));
 sky130_fd_sc_hd__and2_1 _16343_ (.A(_07467_),
    .B(_07479_),
    .X(_07480_));
 sky130_fd_sc_hd__nor2_1 _16344_ (.A(_07467_),
    .B(_07479_),
    .Y(_07481_));
 sky130_fd_sc_hd__or2_1 _16345_ (.A(_07480_),
    .B(_07481_),
    .X(_07482_));
 sky130_fd_sc_hd__o21ba_1 _16346_ (.A1(_07368_),
    .A2(_07382_),
    .B1_N(_07482_),
    .X(_07483_));
 sky130_fd_sc_hd__or3b_4 _16347_ (.A(_07368_),
    .B(_07382_),
    .C_N(_07482_),
    .X(_07484_));
 sky130_fd_sc_hd__nand2b_4 _16348_ (.A_N(_07483_),
    .B(_07484_),
    .Y(_07485_));
 sky130_fd_sc_hd__a21bo_1 _16349_ (.A1(_07394_),
    .A2(_07395_),
    .B1_N(_07397_),
    .X(_07486_));
 sky130_fd_sc_hd__a21o_2 _16350_ (.A1(_07371_),
    .A2(_07380_),
    .B1(_07377_),
    .X(_07488_));
 sky130_fd_sc_hd__nor2_2 _16351_ (.A(net189),
    .B(_06828_),
    .Y(_07489_));
 sky130_fd_sc_hd__and3_1 _16352_ (.A(net194),
    .B(net173),
    .C(_07489_),
    .X(_07490_));
 sky130_fd_sc_hd__o22a_1 _16353_ (.A1(net189),
    .A2(_06733_),
    .B1(_06828_),
    .B2(_06305_),
    .X(_07491_));
 sky130_fd_sc_hd__nor2_1 _16354_ (.A(_07490_),
    .B(_07491_),
    .Y(_07492_));
 sky130_fd_sc_hd__nand2_1 _16355_ (.A(net137),
    .B(_06935_),
    .Y(_07493_));
 sky130_fd_sc_hd__xnor2_1 _16356_ (.A(_07492_),
    .B(_07493_),
    .Y(_07494_));
 sky130_fd_sc_hd__o21ai_1 _16357_ (.A1(_07388_),
    .A2(_07392_),
    .B1(_07494_),
    .Y(_07495_));
 sky130_fd_sc_hd__or3_1 _16358_ (.A(_07388_),
    .B(_07392_),
    .C(_07494_),
    .X(_07496_));
 sky130_fd_sc_hd__and2_2 _16359_ (.A(_07495_),
    .B(_07496_),
    .X(_07497_));
 sky130_fd_sc_hd__nand2b_1 _16360_ (.A_N(_07049_),
    .B(_07497_),
    .Y(_07499_));
 sky130_fd_sc_hd__xnor2_4 _16361_ (.A(_07049_),
    .B(_07497_),
    .Y(_07500_));
 sky130_fd_sc_hd__xnor2_1 _16362_ (.A(_07488_),
    .B(_07500_),
    .Y(_07501_));
 sky130_fd_sc_hd__and2b_2 _16363_ (.A_N(_07501_),
    .B(_07486_),
    .X(_07502_));
 sky130_fd_sc_hd__and2b_1 _16364_ (.A_N(_07486_),
    .B(_07501_),
    .X(_07503_));
 sky130_fd_sc_hd__or2_4 _16365_ (.A(_07502_),
    .B(_07503_),
    .X(_07504_));
 sky130_fd_sc_hd__nor2_1 _16366_ (.A(_07485_),
    .B(_07504_),
    .Y(_07505_));
 sky130_fd_sc_hd__xor2_4 _16367_ (.A(_07485_),
    .B(_07504_),
    .X(_07506_));
 sky130_fd_sc_hd__a21o_2 _16368_ (.A1(_07386_),
    .A2(_07403_),
    .B1(_07385_),
    .X(_07507_));
 sky130_fd_sc_hd__xor2_4 _16369_ (.A(_07506_),
    .B(_07507_),
    .X(_07508_));
 sky130_fd_sc_hd__o21ba_2 _16370_ (.A1(_07387_),
    .A2(_07401_),
    .B1_N(_07399_),
    .X(_07510_));
 sky130_fd_sc_hd__nand2b_1 _16371_ (.A_N(_07510_),
    .B(_07508_),
    .Y(_07511_));
 sky130_fd_sc_hd__xnor2_4 _16372_ (.A(_07508_),
    .B(_07510_),
    .Y(_07512_));
 sky130_fd_sc_hd__o21a_2 _16373_ (.A1(_07408_),
    .A2(_07414_),
    .B1(_07406_),
    .X(_07513_));
 sky130_fd_sc_hd__nand2b_1 _16374_ (.A_N(_07513_),
    .B(_07512_),
    .Y(_07514_));
 sky130_fd_sc_hd__xnor2_4 _16375_ (.A(_07512_),
    .B(_07513_),
    .Y(_07515_));
 sky130_fd_sc_hd__o21ba_2 _16376_ (.A1(_07410_),
    .A2(_07413_),
    .B1_N(_07409_),
    .X(_07516_));
 sky130_fd_sc_hd__nand2b_1 _16377_ (.A_N(_07516_),
    .B(_07515_),
    .Y(_07517_));
 sky130_fd_sc_hd__xnor2_4 _16378_ (.A(_07515_),
    .B(_07516_),
    .Y(_07518_));
 sky130_fd_sc_hd__a21bo_2 _16379_ (.A1(_07415_),
    .A2(_07416_),
    .B1_N(_07419_),
    .X(_07519_));
 sky130_fd_sc_hd__nand2_1 _16380_ (.A(_07518_),
    .B(_07519_),
    .Y(_07521_));
 sky130_fd_sc_hd__xor2_4 _16381_ (.A(_07518_),
    .B(_07519_),
    .X(_07522_));
 sky130_fd_sc_hd__or2_1 _16382_ (.A(_07323_),
    .B(_07421_),
    .X(_07523_));
 sky130_fd_sc_hd__o21a_2 _16383_ (.A1(_07327_),
    .A2(_07523_),
    .B1(_07423_),
    .X(_07524_));
 sky130_fd_sc_hd__nand2_1 _16384_ (.A(_07522_),
    .B(_07524_),
    .Y(_07525_));
 sky130_fd_sc_hd__xor2_4 _16385_ (.A(_07522_),
    .B(_07524_),
    .X(_07526_));
 sky130_fd_sc_hd__nand2_1 _16386_ (.A(net281),
    .B(_07526_),
    .Y(_07527_));
 sky130_fd_sc_hd__or3_2 _16387_ (.A(_01996_),
    .B(_02510_),
    .C(_02511_),
    .X(_07528_));
 sky130_fd_sc_hd__o21ai_4 _16388_ (.A1(_02510_),
    .A2(_02511_),
    .B1(_01996_),
    .Y(_07529_));
 sky130_fd_sc_hd__nand3_4 _16389_ (.A(net261),
    .B(_07528_),
    .C(_07529_),
    .Y(_07530_));
 sky130_fd_sc_hd__a21boi_4 _16390_ (.A1(net424),
    .A2(net274),
    .B1_N(net735),
    .Y(_07532_));
 sky130_fd_sc_hd__nor2_1 _16391_ (.A(net735),
    .B(net271),
    .Y(_07533_));
 sky130_fd_sc_hd__a21o_1 _16392_ (.A1(net424),
    .A2(_07533_),
    .B1(_07532_),
    .X(_07534_));
 sky130_fd_sc_hd__o21ai_2 _16393_ (.A1(_07333_),
    .A2(_07337_),
    .B1(_07431_),
    .Y(_07535_));
 sky130_fd_sc_hd__and2_1 _16394_ (.A(_07430_),
    .B(_07535_),
    .X(_07536_));
 sky130_fd_sc_hd__a21oi_2 _16395_ (.A1(_07430_),
    .A2(_07535_),
    .B1(_07534_),
    .Y(_07537_));
 sky130_fd_sc_hd__xnor2_1 _16396_ (.A(_07534_),
    .B(_07536_),
    .Y(_07538_));
 sky130_fd_sc_hd__nand2b_1 _16397_ (.A_N(_03025_),
    .B(_05775_),
    .Y(_07539_));
 sky130_fd_sc_hd__xor2_1 _16398_ (.A(_05818_),
    .B(_07539_),
    .X(_07540_));
 sky130_fd_sc_hd__nor2_1 _16399_ (.A(net735),
    .B(_05866_),
    .Y(_07541_));
 sky130_fd_sc_hd__or3_1 _16400_ (.A(net251),
    .B(_05868_),
    .C(_07541_),
    .X(_07543_));
 sky130_fd_sc_hd__a221o_1 _16401_ (.A1(_05775_),
    .A2(net239),
    .B1(net232),
    .B2(net735),
    .C1(net245),
    .X(_07544_));
 sky130_fd_sc_hd__a21oi_1 _16402_ (.A1(_03025_),
    .A2(net236),
    .B1(_07544_),
    .Y(_07545_));
 sky130_fd_sc_hd__o22a_1 _16403_ (.A1(net210),
    .A2(_04975_),
    .B1(net202),
    .B2(_06063_),
    .X(_07546_));
 sky130_fd_sc_hd__and3_1 _16404_ (.A(_07543_),
    .B(_07545_),
    .C(_07546_),
    .X(_07547_));
 sky130_fd_sc_hd__o221a_1 _16405_ (.A1(net229),
    .A2(_07538_),
    .B1(_07540_),
    .B2(net253),
    .C1(_07547_),
    .X(_07548_));
 sky130_fd_sc_hd__a32o_1 _16406_ (.A1(_07527_),
    .A2(_07530_),
    .A3(_07548_),
    .B1(net247),
    .B2(net736),
    .X(_07549_));
 sky130_fd_sc_hd__inv_2 _16407_ (.A(_07549_),
    .Y(_08693_));
 sky130_fd_sc_hd__a22o_1 _16408_ (.A1(net452),
    .A2(net199),
    .B1(net197),
    .B2(_07008_),
    .X(_07550_));
 sky130_fd_sc_hd__nor2_1 _16409_ (.A(net196),
    .B(_07129_),
    .Y(_07551_));
 sky130_fd_sc_hd__or3_1 _16410_ (.A(net196),
    .B(net168),
    .C(_07451_),
    .X(_07553_));
 sky130_fd_sc_hd__and2_2 _16411_ (.A(_07550_),
    .B(_07553_),
    .X(_07554_));
 sky130_fd_sc_hd__o21ai_4 _16412_ (.A1(_07450_),
    .A2(_07451_),
    .B1(_07449_),
    .Y(_07555_));
 sky130_fd_sc_hd__nand2_2 _16413_ (.A(_07554_),
    .B(_07555_),
    .Y(_07556_));
 sky130_fd_sc_hd__xor2_2 _16414_ (.A(_07554_),
    .B(_07555_),
    .X(_07557_));
 sky130_fd_sc_hd__a2bb2o_1 _16415_ (.A1_N(net133),
    .A2_N(net171),
    .B1(_06906_),
    .B2(_06313_),
    .X(_07558_));
 sky130_fd_sc_hd__or4_4 _16416_ (.A(net191),
    .B(net133),
    .C(net171),
    .D(net169),
    .X(_07559_));
 sky130_fd_sc_hd__nand2_1 _16417_ (.A(_07558_),
    .B(_07559_),
    .Y(_07560_));
 sky130_fd_sc_hd__or2_2 _16418_ (.A(_06714_),
    .B(_07560_),
    .X(_07561_));
 sky130_fd_sc_hd__xnor2_1 _16419_ (.A(_06714_),
    .B(_07560_),
    .Y(_07562_));
 sky130_fd_sc_hd__inv_2 _16420_ (.A(_07562_),
    .Y(_07564_));
 sky130_fd_sc_hd__or2_1 _16421_ (.A(_07557_),
    .B(_07564_),
    .X(_07565_));
 sky130_fd_sc_hd__nand2_2 _16422_ (.A(_07557_),
    .B(_07564_),
    .Y(_07566_));
 sky130_fd_sc_hd__nand2_1 _16423_ (.A(_07565_),
    .B(_07566_),
    .Y(_07567_));
 sky130_fd_sc_hd__o211a_2 _16424_ (.A1(_07455_),
    .A2(_07463_),
    .B1(_07565_),
    .C1(_07566_),
    .X(_07568_));
 sky130_fd_sc_hd__or3b_2 _16425_ (.A(_07455_),
    .B(_07463_),
    .C_N(_07567_),
    .X(_07569_));
 sky130_fd_sc_hd__nand2b_2 _16426_ (.A_N(_07568_),
    .B(_07569_),
    .Y(_07570_));
 sky130_fd_sc_hd__o21ai_4 _16427_ (.A1(_07469_),
    .A2(_07472_),
    .B1(_07470_),
    .Y(_07571_));
 sky130_fd_sc_hd__a21bo_4 _16428_ (.A1(_07457_),
    .A2(_07460_),
    .B1_N(_07458_),
    .X(_07572_));
 sky130_fd_sc_hd__o22a_1 _16429_ (.A1(net183),
    .A2(net179),
    .B1(net175),
    .B2(net185),
    .X(_07573_));
 sky130_fd_sc_hd__and4_1 _16430_ (.A(_06530_),
    .B(net184),
    .C(net182),
    .D(net177),
    .X(_07575_));
 sky130_fd_sc_hd__nor2_1 _16431_ (.A(_07573_),
    .B(_07575_),
    .Y(_07576_));
 sky130_fd_sc_hd__and3_1 _16432_ (.A(net132),
    .B(net173),
    .C(_07576_),
    .X(_07577_));
 sky130_fd_sc_hd__a21oi_1 _16433_ (.A1(net132),
    .A2(net173),
    .B1(_07576_),
    .Y(_07578_));
 sky130_fd_sc_hd__or2_4 _16434_ (.A(_07577_),
    .B(_07578_),
    .X(_07579_));
 sky130_fd_sc_hd__and2b_1 _16435_ (.A_N(_07579_),
    .B(_07572_),
    .X(_07580_));
 sky130_fd_sc_hd__xnor2_4 _16436_ (.A(_07572_),
    .B(_07579_),
    .Y(_07581_));
 sky130_fd_sc_hd__xnor2_4 _16437_ (.A(_07571_),
    .B(_07581_),
    .Y(_07582_));
 sky130_fd_sc_hd__nor2_2 _16438_ (.A(_07570_),
    .B(_07582_),
    .Y(_07583_));
 sky130_fd_sc_hd__xor2_2 _16439_ (.A(_07570_),
    .B(_07582_),
    .X(_07584_));
 sky130_fd_sc_hd__a21o_1 _16440_ (.A1(_07464_),
    .A2(_07466_),
    .B1(_07480_),
    .X(_07586_));
 sky130_fd_sc_hd__nand2_1 _16441_ (.A(_07584_),
    .B(_07586_),
    .Y(_07587_));
 sky130_fd_sc_hd__xor2_1 _16442_ (.A(_07584_),
    .B(_07586_),
    .X(_07588_));
 sky130_fd_sc_hd__nand2_1 _16443_ (.A(_07495_),
    .B(_07499_),
    .Y(_07589_));
 sky130_fd_sc_hd__or2_2 _16444_ (.A(_07474_),
    .B(_07478_),
    .X(_07590_));
 sky130_fd_sc_hd__nor2_1 _16445_ (.A(net189),
    .B(_06936_),
    .Y(_07591_));
 sky130_fd_sc_hd__or4_2 _16446_ (.A(_06305_),
    .B(net189),
    .C(_06828_),
    .D(_06936_),
    .X(_07592_));
 sky130_fd_sc_hd__a21oi_4 _16447_ (.A1(net195),
    .A2(_06935_),
    .B1(_07489_),
    .Y(_07593_));
 sky130_fd_sc_hd__a31o_2 _16448_ (.A1(net195),
    .A2(_06827_),
    .A3(_07591_),
    .B1(_07593_),
    .X(_07594_));
 sky130_fd_sc_hd__nand2_4 _16449_ (.A(net137),
    .B(_07047_),
    .Y(_07595_));
 sky130_fd_sc_hd__xor2_4 _16450_ (.A(_07594_),
    .B(_07595_),
    .X(_07597_));
 sky130_fd_sc_hd__o21ba_1 _16451_ (.A1(_07491_),
    .A2(_07493_),
    .B1_N(_07490_),
    .X(_07598_));
 sky130_fd_sc_hd__nand2b_1 _16452_ (.A_N(_07598_),
    .B(_07597_),
    .Y(_07599_));
 sky130_fd_sc_hd__xnor2_2 _16453_ (.A(_07597_),
    .B(_07598_),
    .Y(_07600_));
 sky130_fd_sc_hd__xor2_2 _16454_ (.A(_07166_),
    .B(_07600_),
    .X(_07601_));
 sky130_fd_sc_hd__xnor2_1 _16455_ (.A(_07590_),
    .B(_07601_),
    .Y(_07602_));
 sky130_fd_sc_hd__nand2b_1 _16456_ (.A_N(_07602_),
    .B(_07589_),
    .Y(_07603_));
 sky130_fd_sc_hd__xnor2_1 _16457_ (.A(_07589_),
    .B(_07602_),
    .Y(_07604_));
 sky130_fd_sc_hd__nand2_1 _16458_ (.A(_07588_),
    .B(_07604_),
    .Y(_07605_));
 sky130_fd_sc_hd__or2_1 _16459_ (.A(_07588_),
    .B(_07604_),
    .X(_07606_));
 sky130_fd_sc_hd__nand2_1 _16460_ (.A(_07605_),
    .B(_07606_),
    .Y(_07608_));
 sky130_fd_sc_hd__o21ba_1 _16461_ (.A1(_07483_),
    .A2(_07505_),
    .B1_N(_07608_),
    .X(_07609_));
 sky130_fd_sc_hd__or3b_2 _16462_ (.A(_07483_),
    .B(_07505_),
    .C_N(_07608_),
    .X(_07610_));
 sky130_fd_sc_hd__nand2b_4 _16463_ (.A_N(_07609_),
    .B(_07610_),
    .Y(_07611_));
 sky130_fd_sc_hd__a21oi_4 _16464_ (.A1(_07488_),
    .A2(_07500_),
    .B1(_07502_),
    .Y(_07612_));
 sky130_fd_sc_hd__nor2_1 _16465_ (.A(_07611_),
    .B(_07612_),
    .Y(_07613_));
 sky130_fd_sc_hd__xnor2_4 _16466_ (.A(_07611_),
    .B(_07612_),
    .Y(_07614_));
 sky130_fd_sc_hd__a21bo_2 _16467_ (.A1(_07506_),
    .A2(_07507_),
    .B1_N(_07511_),
    .X(_07615_));
 sky130_fd_sc_hd__and2b_2 _16468_ (.A_N(_07614_),
    .B(_07615_),
    .X(_07616_));
 sky130_fd_sc_hd__xor2_4 _16469_ (.A(_07614_),
    .B(_07615_),
    .X(_07617_));
 sky130_fd_sc_hd__and3_1 _16470_ (.A(_07514_),
    .B(_07517_),
    .C(_07617_),
    .X(_07619_));
 sky130_fd_sc_hd__a21oi_2 _16471_ (.A1(_07514_),
    .A2(_07517_),
    .B1(_07617_),
    .Y(_07620_));
 sky130_fd_sc_hd__or2_1 _16472_ (.A(_07619_),
    .B(_07620_),
    .X(_07621_));
 sky130_fd_sc_hd__a21oi_1 _16473_ (.A1(_07521_),
    .A2(_07525_),
    .B1(_07621_),
    .Y(_07622_));
 sky130_fd_sc_hd__a31o_1 _16474_ (.A1(_07521_),
    .A2(_07525_),
    .A3(_07621_),
    .B1(net279),
    .X(_07623_));
 sky130_fd_sc_hd__or2_4 _16475_ (.A(_07622_),
    .B(_07623_),
    .X(_07624_));
 sky130_fd_sc_hd__a21oi_1 _16476_ (.A1(_01995_),
    .A2(_07529_),
    .B1(_02024_),
    .Y(_07625_));
 sky130_fd_sc_hd__a31o_1 _16477_ (.A1(_01995_),
    .A2(_02024_),
    .A3(_07529_),
    .B1(net256),
    .X(_07626_));
 sky130_fd_sc_hd__or2_4 _16478_ (.A(_07625_),
    .B(_07626_),
    .X(_07627_));
 sky130_fd_sc_hd__a21bo_1 _16479_ (.A1(net415),
    .A2(net274),
    .B1_N(net727),
    .X(_07628_));
 sky130_fd_sc_hd__or3b_1 _16480_ (.A(net727),
    .B(net271),
    .C_N(net415),
    .X(_07630_));
 sky130_fd_sc_hd__and2_1 _16481_ (.A(_07628_),
    .B(_07630_),
    .X(_07631_));
 sky130_fd_sc_hd__o21ai_2 _16482_ (.A1(_07532_),
    .A2(_07537_),
    .B1(_07631_),
    .Y(_07632_));
 sky130_fd_sc_hd__o311a_1 _16483_ (.A1(_07532_),
    .A2(_07537_),
    .A3(_07631_),
    .B1(_07632_),
    .C1(net230),
    .X(_07633_));
 sky130_fd_sc_hd__a21o_1 _16484_ (.A1(_03363_),
    .A2(_05774_),
    .B1(_05819_),
    .X(_07634_));
 sky130_fd_sc_hd__nand2_1 _16485_ (.A(net254),
    .B(_07634_),
    .Y(_07635_));
 sky130_fd_sc_hd__a31o_1 _16486_ (.A1(_03363_),
    .A2(_05774_),
    .A3(_05819_),
    .B1(_07635_),
    .X(_07636_));
 sky130_fd_sc_hd__a21oi_1 _16487_ (.A1(net727),
    .A2(_05868_),
    .B1(net251),
    .Y(_07637_));
 sky130_fd_sc_hd__o21ai_1 _16488_ (.A1(net727),
    .A2(_05868_),
    .B1(_07637_),
    .Y(_07638_));
 sky130_fd_sc_hd__a221o_1 _16489_ (.A1(_05774_),
    .A2(net239),
    .B1(net232),
    .B2(net727),
    .C1(net245),
    .X(_07639_));
 sky130_fd_sc_hd__o21ba_1 _16490_ (.A1(_03363_),
    .A2(net235),
    .B1_N(_07639_),
    .X(_07641_));
 sky130_fd_sc_hd__o22a_1 _16491_ (.A1(net210),
    .A2(_05074_),
    .B1(net202),
    .B2(_06132_),
    .X(_07642_));
 sky130_fd_sc_hd__and3_1 _16492_ (.A(_07638_),
    .B(_07641_),
    .C(_07642_),
    .X(_07643_));
 sky130_fd_sc_hd__and3b_1 _16493_ (.A_N(_07633_),
    .B(_07636_),
    .C(_07643_),
    .X(_07644_));
 sky130_fd_sc_hd__a32o_1 _16494_ (.A1(_07624_),
    .A2(_07627_),
    .A3(_07644_),
    .B1(net247),
    .B2(net728),
    .X(_07645_));
 sky130_fd_sc_hd__inv_2 _16495_ (.A(_07645_),
    .Y(_08694_));
 sky130_fd_sc_hd__o22ai_1 _16496_ (.A1(net187),
    .A2(net171),
    .B1(net169),
    .B2(net133),
    .Y(_07646_));
 sky130_fd_sc_hd__or4_2 _16497_ (.A(net133),
    .B(net187),
    .C(net171),
    .D(net169),
    .X(_07647_));
 sky130_fd_sc_hd__nand2_1 _16498_ (.A(_07646_),
    .B(_07647_),
    .Y(_07648_));
 sky130_fd_sc_hd__or3_2 _16499_ (.A(net183),
    .B(_06712_),
    .C(_07648_),
    .X(_07649_));
 sky130_fd_sc_hd__o21ai_1 _16500_ (.A1(net183),
    .A2(_06712_),
    .B1(_07648_),
    .Y(_07651_));
 sky130_fd_sc_hd__and2_2 _16501_ (.A(_07649_),
    .B(_07651_),
    .X(_07652_));
 sky130_fd_sc_hd__nor2_2 _16502_ (.A(net191),
    .B(_07009_),
    .Y(_07653_));
 sky130_fd_sc_hd__nand2_1 _16503_ (.A(_07551_),
    .B(_07653_),
    .Y(_07654_));
 sky130_fd_sc_hd__nand2b_1 _16504_ (.A_N(_07654_),
    .B(_07451_),
    .Y(_07655_));
 sky130_fd_sc_hd__or2_1 _16505_ (.A(_06313_),
    .B(_07553_),
    .X(_07656_));
 sky130_fd_sc_hd__o211a_2 _16506_ (.A1(_07551_),
    .A2(_07653_),
    .B1(_07655_),
    .C1(_07656_),
    .X(_07657_));
 sky130_fd_sc_hd__xnor2_2 _16507_ (.A(_07652_),
    .B(_07657_),
    .Y(_07658_));
 sky130_fd_sc_hd__a21oi_4 _16508_ (.A1(_07556_),
    .A2(_07566_),
    .B1(_07658_),
    .Y(_07659_));
 sky130_fd_sc_hd__and3_1 _16509_ (.A(_07556_),
    .B(_07566_),
    .C(_07658_),
    .X(_07660_));
 sky130_fd_sc_hd__or2_1 _16510_ (.A(_07659_),
    .B(_07660_),
    .X(_07662_));
 sky130_fd_sc_hd__or2_1 _16511_ (.A(_07575_),
    .B(_07577_),
    .X(_07663_));
 sky130_fd_sc_hd__nand2_1 _16512_ (.A(_06530_),
    .B(net173),
    .Y(_07664_));
 sky130_fd_sc_hd__o21ai_1 _16513_ (.A1(net179),
    .A2(net175),
    .B1(_07664_),
    .Y(_07665_));
 sky130_fd_sc_hd__or3_2 _16514_ (.A(net179),
    .B(net175),
    .C(_07664_),
    .X(_07666_));
 sky130_fd_sc_hd__nand2_2 _16515_ (.A(_07665_),
    .B(_07666_),
    .Y(_07667_));
 sky130_fd_sc_hd__nand2_2 _16516_ (.A(net797),
    .B(net132),
    .Y(_07668_));
 sky130_fd_sc_hd__xnor2_2 _16517_ (.A(_07667_),
    .B(_07668_),
    .Y(_07669_));
 sky130_fd_sc_hd__a21oi_2 _16518_ (.A1(_07559_),
    .A2(_07561_),
    .B1(_07669_),
    .Y(_07670_));
 sky130_fd_sc_hd__and3_1 _16519_ (.A(_07559_),
    .B(_07561_),
    .C(_07669_),
    .X(_07671_));
 sky130_fd_sc_hd__nor2_1 _16520_ (.A(_07670_),
    .B(_07671_),
    .Y(_07673_));
 sky130_fd_sc_hd__and2_1 _16521_ (.A(_07663_),
    .B(_07673_),
    .X(_07674_));
 sky130_fd_sc_hd__xnor2_1 _16522_ (.A(_07663_),
    .B(_07673_),
    .Y(_07675_));
 sky130_fd_sc_hd__nor2_2 _16523_ (.A(_07662_),
    .B(_07675_),
    .Y(_07676_));
 sky130_fd_sc_hd__and2_1 _16524_ (.A(_07662_),
    .B(_07675_),
    .X(_07677_));
 sky130_fd_sc_hd__nor2_2 _16525_ (.A(_07676_),
    .B(_07677_),
    .Y(_07678_));
 sky130_fd_sc_hd__o21ai_4 _16526_ (.A1(_07568_),
    .A2(_07583_),
    .B1(_07678_),
    .Y(_07679_));
 sky130_fd_sc_hd__or3_1 _16527_ (.A(_07568_),
    .B(_07583_),
    .C(_07678_),
    .X(_07680_));
 sky130_fd_sc_hd__and2_1 _16528_ (.A(_07679_),
    .B(_07680_),
    .X(_07681_));
 sky130_fd_sc_hd__a21bo_1 _16529_ (.A1(_07166_),
    .A2(_07600_),
    .B1_N(_07599_),
    .X(_07682_));
 sky130_fd_sc_hd__a21o_1 _16530_ (.A1(_07571_),
    .A2(_07581_),
    .B1(_07580_),
    .X(_07684_));
 sky130_fd_sc_hd__nand2_1 _16531_ (.A(net195),
    .B(_07047_),
    .Y(_07685_));
 sky130_fd_sc_hd__and2b_1 _16532_ (.A_N(_07591_),
    .B(_07685_),
    .X(_07686_));
 sky130_fd_sc_hd__and3_2 _16533_ (.A(net195),
    .B(_07047_),
    .C(_07591_),
    .X(_07687_));
 sky130_fd_sc_hd__nor2_4 _16534_ (.A(_07686_),
    .B(_07687_),
    .Y(_07688_));
 sky130_fd_sc_hd__nand2_2 _16535_ (.A(net137),
    .B(_07164_),
    .Y(_07689_));
 sky130_fd_sc_hd__and3_1 _16536_ (.A(net137),
    .B(_07164_),
    .C(_07688_),
    .X(_07690_));
 sky130_fd_sc_hd__xnor2_4 _16537_ (.A(_07688_),
    .B(_07689_),
    .Y(_07691_));
 sky130_fd_sc_hd__o21ai_4 _16538_ (.A1(_07593_),
    .A2(_07595_),
    .B1(_07592_),
    .Y(_07692_));
 sky130_fd_sc_hd__nand2_4 _16539_ (.A(_07691_),
    .B(_07692_),
    .Y(_07693_));
 sky130_fd_sc_hd__inv_2 _16540_ (.A(_07693_),
    .Y(_07695_));
 sky130_fd_sc_hd__nor2_1 _16541_ (.A(_07691_),
    .B(_07692_),
    .Y(_07696_));
 sky130_fd_sc_hd__nor2_2 _16542_ (.A(_07695_),
    .B(_07696_),
    .Y(_07697_));
 sky130_fd_sc_hd__xnor2_1 _16543_ (.A(_07684_),
    .B(_07697_),
    .Y(_07698_));
 sky130_fd_sc_hd__and2b_1 _16544_ (.A_N(_07698_),
    .B(_07682_),
    .X(_07699_));
 sky130_fd_sc_hd__xnor2_1 _16545_ (.A(_07682_),
    .B(_07698_),
    .Y(_07700_));
 sky130_fd_sc_hd__nand2_2 _16546_ (.A(_07681_),
    .B(_07700_),
    .Y(_07701_));
 sky130_fd_sc_hd__or2_1 _16547_ (.A(_07681_),
    .B(_07700_),
    .X(_07702_));
 sky130_fd_sc_hd__nand2_1 _16548_ (.A(_07701_),
    .B(_07702_),
    .Y(_07703_));
 sky130_fd_sc_hd__a21o_2 _16549_ (.A1(_07587_),
    .A2(_07605_),
    .B1(_07703_),
    .X(_07704_));
 sky130_fd_sc_hd__nand3_1 _16550_ (.A(_07587_),
    .B(_07605_),
    .C(_07703_),
    .Y(_07706_));
 sky130_fd_sc_hd__nand2_2 _16551_ (.A(_07704_),
    .B(_07706_),
    .Y(_07707_));
 sky130_fd_sc_hd__a21bo_2 _16552_ (.A1(_07590_),
    .A2(_07601_),
    .B1_N(_07603_),
    .X(_07708_));
 sky130_fd_sc_hd__nand2b_2 _16553_ (.A_N(_07707_),
    .B(_07708_),
    .Y(_07709_));
 sky130_fd_sc_hd__xnor2_2 _16554_ (.A(_07707_),
    .B(_07708_),
    .Y(_07710_));
 sky130_fd_sc_hd__o21a_4 _16555_ (.A1(_07609_),
    .A2(_07613_),
    .B1(_07710_),
    .X(_07711_));
 sky130_fd_sc_hd__inv_2 _16556_ (.A(_07711_),
    .Y(_07712_));
 sky130_fd_sc_hd__or3_4 _16557_ (.A(_07609_),
    .B(_07613_),
    .C(_07710_),
    .X(_07713_));
 sky130_fd_sc_hd__nand3_4 _16558_ (.A(_07616_),
    .B(_07712_),
    .C(_07713_),
    .Y(_07714_));
 sky130_fd_sc_hd__a21o_1 _16559_ (.A1(_07712_),
    .A2(_07713_),
    .B1(_07616_),
    .X(_07715_));
 sky130_fd_sc_hd__nand2_2 _16560_ (.A(_07714_),
    .B(_07715_),
    .Y(_07717_));
 sky130_fd_sc_hd__or3b_2 _16561_ (.A(_07619_),
    .B(_07620_),
    .C_N(_07522_),
    .X(_07718_));
 sky130_fd_sc_hd__nand3b_1 _16562_ (.A_N(_07718_),
    .B(_07523_),
    .C(_07423_),
    .Y(_07719_));
 sky130_fd_sc_hd__nor2_1 _16563_ (.A(_07521_),
    .B(_07619_),
    .Y(_07720_));
 sky130_fd_sc_hd__nor2_1 _16564_ (.A(_07620_),
    .B(_07720_),
    .Y(_07721_));
 sky130_fd_sc_hd__o311a_4 _16565_ (.A1(_07328_),
    .A2(_07424_),
    .A3(_07718_),
    .B1(_07719_),
    .C1(_07721_),
    .X(_07722_));
 sky130_fd_sc_hd__nor2_2 _16566_ (.A(_07717_),
    .B(_07722_),
    .Y(_07723_));
 sky130_fd_sc_hd__a21o_1 _16567_ (.A1(_07717_),
    .A2(_07722_),
    .B1(net278),
    .X(_07724_));
 sky130_fd_sc_hd__nor2_1 _16568_ (.A(_02513_),
    .B(_02551_),
    .Y(_07725_));
 sky130_fd_sc_hd__a211o_4 _16569_ (.A1(_02513_),
    .A2(_02551_),
    .B1(net256),
    .C1(_07725_),
    .X(_07726_));
 sky130_fd_sc_hd__a21bo_1 _16570_ (.A1(net409),
    .A2(net274),
    .B1_N(net718),
    .X(_07728_));
 sky130_fd_sc_hd__or3b_1 _16571_ (.A(net717),
    .B(net271),
    .C_N(net409),
    .X(_07729_));
 sky130_fd_sc_hd__nand2_1 _16572_ (.A(_07728_),
    .B(_07729_),
    .Y(_07730_));
 sky130_fd_sc_hd__a21o_1 _16573_ (.A1(_07628_),
    .A2(_07632_),
    .B1(_07730_),
    .X(_07731_));
 sky130_fd_sc_hd__nand2_1 _16574_ (.A(net230),
    .B(_07731_),
    .Y(_07732_));
 sky130_fd_sc_hd__a31o_1 _16575_ (.A1(_07628_),
    .A2(_07632_),
    .A3(_07730_),
    .B1(_07732_),
    .X(_07733_));
 sky130_fd_sc_hd__nand2b_1 _16576_ (.A_N(_03365_),
    .B(_05773_),
    .Y(_07734_));
 sky130_fd_sc_hd__xor2_1 _16577_ (.A(_05820_),
    .B(_07734_),
    .X(_07735_));
 sky130_fd_sc_hd__a21oi_1 _16578_ (.A1(net727),
    .A2(_05868_),
    .B1(net717),
    .Y(_07736_));
 sky130_fd_sc_hd__or3_2 _16579_ (.A(net251),
    .B(_05869_),
    .C(_07736_),
    .X(_07737_));
 sky130_fd_sc_hd__a221o_1 _16580_ (.A1(_05773_),
    .A2(net239),
    .B1(net233),
    .B2(net717),
    .C1(net245),
    .X(_07739_));
 sky130_fd_sc_hd__a21oi_1 _16581_ (.A1(_03365_),
    .A2(net236),
    .B1(_07739_),
    .Y(_07740_));
 sky130_fd_sc_hd__or2_1 _16582_ (.A(net202),
    .B(_06216_),
    .X(_07741_));
 sky130_fd_sc_hd__o211a_1 _16583_ (.A1(net211),
    .A2(_05163_),
    .B1(_07740_),
    .C1(_07741_),
    .X(_07742_));
 sky130_fd_sc_hd__o211a_1 _16584_ (.A1(net252),
    .A2(_07735_),
    .B1(_07742_),
    .C1(_07726_),
    .X(_07743_));
 sky130_fd_sc_hd__o211a_1 _16585_ (.A1(_07723_),
    .A2(_07724_),
    .B1(_07737_),
    .C1(_07743_),
    .X(_07744_));
 sky130_fd_sc_hd__a22oi_4 _16586_ (.A1(net718),
    .A2(net247),
    .B1(_07733_),
    .B2(_07744_),
    .Y(_08696_));
 sky130_fd_sc_hd__o21ai_1 _16587_ (.A1(_07717_),
    .A2(_07722_),
    .B1(_07714_),
    .Y(_07745_));
 sky130_fd_sc_hd__o22a_1 _16588_ (.A1(net183),
    .A2(net171),
    .B1(net169),
    .B2(net187),
    .X(_07746_));
 sky130_fd_sc_hd__and4_2 _16589_ (.A(net188),
    .B(net184),
    .C(net172),
    .D(net170),
    .X(_07747_));
 sky130_fd_sc_hd__nor2_1 _16590_ (.A(_07746_),
    .B(_07747_),
    .Y(_07749_));
 sky130_fd_sc_hd__and3_2 _16591_ (.A(net177),
    .B(net223),
    .C(_07749_),
    .X(_07750_));
 sky130_fd_sc_hd__a21oi_1 _16592_ (.A1(net177),
    .A2(net223),
    .B1(_07749_),
    .Y(_07751_));
 sky130_fd_sc_hd__nor2_2 _16593_ (.A(_07750_),
    .B(_07751_),
    .Y(_07752_));
 sky130_fd_sc_hd__nor2_4 _16594_ (.A(net133),
    .B(_07009_),
    .Y(_07753_));
 sky130_fd_sc_hd__or3b_4 _16595_ (.A(net191),
    .B(net168),
    .C_N(_07654_),
    .X(_07754_));
 sky130_fd_sc_hd__xnor2_4 _16596_ (.A(_07753_),
    .B(_07754_),
    .Y(_07755_));
 sky130_fd_sc_hd__xnor2_2 _16597_ (.A(_07752_),
    .B(_07755_),
    .Y(_07756_));
 sky130_fd_sc_hd__a21boi_2 _16598_ (.A1(_07652_),
    .A2(_07657_),
    .B1_N(_07656_),
    .Y(_07757_));
 sky130_fd_sc_hd__nand2_1 _16599_ (.A(_07756_),
    .B(_07757_),
    .Y(_07758_));
 sky130_fd_sc_hd__or2_1 _16600_ (.A(_07756_),
    .B(_07757_),
    .X(_07760_));
 sky130_fd_sc_hd__nand2_1 _16601_ (.A(_07758_),
    .B(_07760_),
    .Y(_07761_));
 sky130_fd_sc_hd__o21ai_1 _16602_ (.A1(_07667_),
    .A2(_07668_),
    .B1(_07666_),
    .Y(_07762_));
 sky130_fd_sc_hd__a22o_1 _16603_ (.A1(net182),
    .A2(net173),
    .B1(_06827_),
    .B2(_06530_),
    .X(_07763_));
 sky130_fd_sc_hd__and4_1 _16604_ (.A(net798),
    .B(_06530_),
    .C(net182),
    .D(net174),
    .X(_07764_));
 sky130_fd_sc_hd__o31a_2 _16605_ (.A1(net179),
    .A2(_06828_),
    .A3(_07664_),
    .B1(_07763_),
    .X(_07765_));
 sky130_fd_sc_hd__nand2_1 _16606_ (.A(net784),
    .B(net132),
    .Y(_07766_));
 sky130_fd_sc_hd__xor2_2 _16607_ (.A(_07765_),
    .B(_07766_),
    .X(_07767_));
 sky130_fd_sc_hd__a21oi_2 _16608_ (.A1(_07647_),
    .A2(_07649_),
    .B1(_07767_),
    .Y(_07768_));
 sky130_fd_sc_hd__and3_1 _16609_ (.A(_07647_),
    .B(_07649_),
    .C(_07767_),
    .X(_07769_));
 sky130_fd_sc_hd__or2_1 _16610_ (.A(_07768_),
    .B(_07769_),
    .X(_07771_));
 sky130_fd_sc_hd__and2b_1 _16611_ (.A_N(_07771_),
    .B(_07762_),
    .X(_07772_));
 sky130_fd_sc_hd__and2b_1 _16612_ (.A_N(_07762_),
    .B(_07771_),
    .X(_07773_));
 sky130_fd_sc_hd__nor2_1 _16613_ (.A(_07772_),
    .B(_07773_),
    .Y(_07774_));
 sky130_fd_sc_hd__xnor2_1 _16614_ (.A(_07761_),
    .B(_07774_),
    .Y(_07775_));
 sky130_fd_sc_hd__o21a_1 _16615_ (.A1(_07659_),
    .A2(_07676_),
    .B1(_07775_),
    .X(_07776_));
 sky130_fd_sc_hd__nor3_1 _16616_ (.A(_07659_),
    .B(_07676_),
    .C(_07775_),
    .Y(_07777_));
 sky130_fd_sc_hd__nor2_2 _16617_ (.A(_07776_),
    .B(_07777_),
    .Y(_07778_));
 sky130_fd_sc_hd__a22o_1 _16618_ (.A1(_06372_),
    .A2(_07047_),
    .B1(_07164_),
    .B2(net195),
    .X(_07779_));
 sky130_fd_sc_hd__or3_4 _16619_ (.A(net189),
    .B(_07165_),
    .C(_07685_),
    .X(_07780_));
 sky130_fd_sc_hd__and2_1 _16620_ (.A(_07779_),
    .B(_07780_),
    .X(_07782_));
 sky130_fd_sc_hd__o21a_1 _16621_ (.A1(_07687_),
    .A2(_07690_),
    .B1(_07782_),
    .X(_07783_));
 sky130_fd_sc_hd__nor3_1 _16622_ (.A(_07687_),
    .B(_07690_),
    .C(_07782_),
    .Y(_07784_));
 sky130_fd_sc_hd__or2_1 _16623_ (.A(_07783_),
    .B(_07784_),
    .X(_07785_));
 sky130_fd_sc_hd__o21ba_2 _16624_ (.A1(_07670_),
    .A2(_07674_),
    .B1_N(_07785_),
    .X(_07786_));
 sky130_fd_sc_hd__or3b_4 _16625_ (.A(_07670_),
    .B(_07674_),
    .C_N(_07785_),
    .X(_07787_));
 sky130_fd_sc_hd__and2b_2 _16626_ (.A_N(_07786_),
    .B(_07787_),
    .X(_07788_));
 sky130_fd_sc_hd__xnor2_4 _16627_ (.A(_07693_),
    .B(_07788_),
    .Y(_07789_));
 sky130_fd_sc_hd__xnor2_2 _16628_ (.A(_07778_),
    .B(_07789_),
    .Y(_07790_));
 sky130_fd_sc_hd__a21oi_4 _16629_ (.A1(_07679_),
    .A2(_07701_),
    .B1(_07790_),
    .Y(_07791_));
 sky130_fd_sc_hd__and3_1 _16630_ (.A(_07679_),
    .B(_07701_),
    .C(_07790_),
    .X(_07793_));
 sky130_fd_sc_hd__or2_2 _16631_ (.A(_07791_),
    .B(_07793_),
    .X(_07794_));
 sky130_fd_sc_hd__a21oi_2 _16632_ (.A1(_07684_),
    .A2(_07697_),
    .B1(_07699_),
    .Y(_07795_));
 sky130_fd_sc_hd__nor2_2 _16633_ (.A(_07794_),
    .B(_07795_),
    .Y(_07796_));
 sky130_fd_sc_hd__xnor2_1 _16634_ (.A(_07794_),
    .B(_07795_),
    .Y(_07797_));
 sky130_fd_sc_hd__a21oi_2 _16635_ (.A1(_07704_),
    .A2(_07709_),
    .B1(_07797_),
    .Y(_07798_));
 sky130_fd_sc_hd__and3_1 _16636_ (.A(_07704_),
    .B(_07709_),
    .C(_07797_),
    .X(_07799_));
 sky130_fd_sc_hd__or2_4 _16637_ (.A(_07798_),
    .B(_07799_),
    .X(_07800_));
 sky130_fd_sc_hd__xnor2_4 _16638_ (.A(_07711_),
    .B(_07800_),
    .Y(_07801_));
 sky130_fd_sc_hd__xnor2_1 _16639_ (.A(_07745_),
    .B(_07801_),
    .Y(_07802_));
 sky130_fd_sc_hd__a22o_2 _16640_ (.A1(_02022_),
    .A2(_02550_),
    .B1(_02551_),
    .B2(_02513_),
    .X(_07804_));
 sky130_fd_sc_hd__xnor2_4 _16641_ (.A(_02554_),
    .B(_07804_),
    .Y(_07805_));
 sky130_fd_sc_hd__a21boi_4 _16642_ (.A1(net402),
    .A2(net275),
    .B1_N(net710),
    .Y(_07806_));
 sky130_fd_sc_hd__inv_2 _16643_ (.A(_07806_),
    .Y(_07807_));
 sky130_fd_sc_hd__and3b_1 _16644_ (.A_N(net710),
    .B(net274),
    .C(net402),
    .X(_07808_));
 sky130_fd_sc_hd__o211a_1 _16645_ (.A1(_07806_),
    .A2(_07808_),
    .B1(_07728_),
    .C1(_07731_),
    .X(_07809_));
 sky130_fd_sc_hd__a211o_1 _16646_ (.A1(_07728_),
    .A2(_07731_),
    .B1(_07806_),
    .C1(_07808_),
    .X(_07810_));
 sky130_fd_sc_hd__inv_2 _16647_ (.A(_07810_),
    .Y(_07811_));
 sky130_fd_sc_hd__or3_1 _16648_ (.A(net229),
    .B(_07809_),
    .C(_07811_),
    .X(_07812_));
 sky130_fd_sc_hd__and3_1 _16649_ (.A(_04070_),
    .B(_05772_),
    .C(_05821_),
    .X(_07813_));
 sky130_fd_sc_hd__a21oi_1 _16650_ (.A1(_04070_),
    .A2(_05772_),
    .B1(_05821_),
    .Y(_07815_));
 sky130_fd_sc_hd__nor2_1 _16651_ (.A(net709),
    .B(_05869_),
    .Y(_07816_));
 sky130_fd_sc_hd__or3_1 _16652_ (.A(net250),
    .B(_05870_),
    .C(_07816_),
    .X(_07817_));
 sky130_fd_sc_hd__or2_1 _16653_ (.A(net208),
    .B(_05247_),
    .X(_07818_));
 sky130_fd_sc_hd__a221o_1 _16654_ (.A1(_05772_),
    .A2(net238),
    .B1(net232),
    .B2(net709),
    .C1(net244),
    .X(_07819_));
 sky130_fd_sc_hd__o21ba_1 _16655_ (.A1(_04070_),
    .A2(net235),
    .B1_N(_07819_),
    .X(_07820_));
 sky130_fd_sc_hd__o211a_1 _16656_ (.A1(net203),
    .A2(_06286_),
    .B1(_07818_),
    .C1(_07820_),
    .X(_07821_));
 sky130_fd_sc_hd__o311a_2 _16657_ (.A1(net252),
    .A2(_07813_),
    .A3(_07815_),
    .B1(_07817_),
    .C1(_07821_),
    .X(_07822_));
 sky130_fd_sc_hd__o211a_1 _16658_ (.A1(net257),
    .A2(_07805_),
    .B1(_07812_),
    .C1(_07822_),
    .X(_07823_));
 sky130_fd_sc_hd__o21a_1 _16659_ (.A1(net278),
    .A2(_07802_),
    .B1(_07823_),
    .X(_07824_));
 sky130_fd_sc_hd__a21oi_4 _16660_ (.A1(net709),
    .A2(net247),
    .B1(_07824_),
    .Y(_08697_));
 sky130_fd_sc_hd__o22a_1 _16661_ (.A1(net175),
    .A2(net171),
    .B1(net169),
    .B2(net183),
    .X(_07826_));
 sky130_fd_sc_hd__or4_2 _16662_ (.A(net183),
    .B(net175),
    .C(net171),
    .D(net169),
    .X(_07827_));
 sky130_fd_sc_hd__nand2b_1 _16663_ (.A_N(_07826_),
    .B(_07827_),
    .Y(_07828_));
 sky130_fd_sc_hd__nand2_1 _16664_ (.A(net223),
    .B(net174),
    .Y(_07829_));
 sky130_fd_sc_hd__xor2_1 _16665_ (.A(_07828_),
    .B(_07829_),
    .X(_07830_));
 sky130_fd_sc_hd__nor2_1 _16666_ (.A(net133),
    .B(net168),
    .Y(_07831_));
 sky130_fd_sc_hd__or4_2 _16667_ (.A(net133),
    .B(net187),
    .C(_07009_),
    .D(net168),
    .X(_07832_));
 sky130_fd_sc_hd__a21oi_1 _16668_ (.A1(_07653_),
    .A2(_07831_),
    .B1(_07832_),
    .Y(_07833_));
 sky130_fd_sc_hd__o32a_1 _16669_ (.A1(net133),
    .A2(net168),
    .A3(_07653_),
    .B1(net187),
    .B2(_07009_),
    .X(_07834_));
 sky130_fd_sc_hd__nand3_2 _16670_ (.A(_07653_),
    .B(_07831_),
    .C(_07832_),
    .Y(_07836_));
 sky130_fd_sc_hd__nor2_1 _16671_ (.A(_07833_),
    .B(_07834_),
    .Y(_07837_));
 sky130_fd_sc_hd__nand2_1 _16672_ (.A(_07830_),
    .B(_07837_),
    .Y(_07838_));
 sky130_fd_sc_hd__or2_1 _16673_ (.A(_07830_),
    .B(_07837_),
    .X(_07839_));
 sky130_fd_sc_hd__nand2_1 _16674_ (.A(_07838_),
    .B(_07839_),
    .Y(_07840_));
 sky130_fd_sc_hd__a2bb2o_1 _16675_ (.A1_N(_07654_),
    .A2_N(_07831_),
    .B1(_07755_),
    .B2(_07752_),
    .X(_07841_));
 sky130_fd_sc_hd__and2b_1 _16676_ (.A_N(_07840_),
    .B(_07841_),
    .X(_07842_));
 sky130_fd_sc_hd__and2b_1 _16677_ (.A_N(_07841_),
    .B(_07840_),
    .X(_07843_));
 sky130_fd_sc_hd__or2_1 _16678_ (.A(_07842_),
    .B(_07843_),
    .X(_07844_));
 sky130_fd_sc_hd__a31o_2 _16679_ (.A1(net785),
    .A2(net132),
    .A3(_07763_),
    .B1(_07764_),
    .X(_07845_));
 sky130_fd_sc_hd__o22a_1 _16680_ (.A1(net179),
    .A2(_06828_),
    .B1(_06936_),
    .B2(net185),
    .X(_07847_));
 sky130_fd_sc_hd__or4_1 _16681_ (.A(net185),
    .B(net179),
    .C(_06828_),
    .D(_06936_),
    .X(_07848_));
 sky130_fd_sc_hd__nand2b_1 _16682_ (.A_N(_07847_),
    .B(_07848_),
    .Y(_07849_));
 sky130_fd_sc_hd__nand2_1 _16683_ (.A(net776),
    .B(net132),
    .Y(_07850_));
 sky130_fd_sc_hd__xnor2_1 _16684_ (.A(_07849_),
    .B(_07850_),
    .Y(_07851_));
 sky130_fd_sc_hd__o21ba_1 _16685_ (.A1(_07747_),
    .A2(_07750_),
    .B1_N(_07851_),
    .X(_07852_));
 sky130_fd_sc_hd__or3b_1 _16686_ (.A(_07747_),
    .B(_07750_),
    .C_N(_07851_),
    .X(_07853_));
 sky130_fd_sc_hd__and2b_1 _16687_ (.A_N(_07852_),
    .B(_07853_),
    .X(_07854_));
 sky130_fd_sc_hd__xor2_2 _16688_ (.A(_07845_),
    .B(_07854_),
    .X(_07855_));
 sky130_fd_sc_hd__and2b_1 _16689_ (.A_N(_07844_),
    .B(_07855_),
    .X(_07856_));
 sky130_fd_sc_hd__xnor2_1 _16690_ (.A(_07844_),
    .B(_07855_),
    .Y(_07858_));
 sky130_fd_sc_hd__a21boi_1 _16691_ (.A1(_07758_),
    .A2(_07774_),
    .B1_N(_07760_),
    .Y(_07859_));
 sky130_fd_sc_hd__nand2b_1 _16692_ (.A_N(_07859_),
    .B(_07858_),
    .Y(_07860_));
 sky130_fd_sc_hd__nand2b_1 _16693_ (.A_N(_07858_),
    .B(_07859_),
    .Y(_07861_));
 sky130_fd_sc_hd__nand2_1 _16694_ (.A(_07860_),
    .B(_07861_),
    .Y(_07862_));
 sky130_fd_sc_hd__and3_1 _16695_ (.A(_06372_),
    .B(_07164_),
    .C(_07685_),
    .X(_07863_));
 sky130_fd_sc_hd__o21ai_1 _16696_ (.A1(_07768_),
    .A2(_07772_),
    .B1(_07863_),
    .Y(_07864_));
 sky130_fd_sc_hd__or3_1 _16697_ (.A(_07768_),
    .B(_07772_),
    .C(_07863_),
    .X(_07865_));
 sky130_fd_sc_hd__and2_1 _16698_ (.A(_07864_),
    .B(_07865_),
    .X(_07866_));
 sky130_fd_sc_hd__xnor2_1 _16699_ (.A(_07783_),
    .B(_07866_),
    .Y(_07867_));
 sky130_fd_sc_hd__or2_2 _16700_ (.A(_07862_),
    .B(_07867_),
    .X(_07869_));
 sky130_fd_sc_hd__nand2_1 _16701_ (.A(_07862_),
    .B(_07867_),
    .Y(_07870_));
 sky130_fd_sc_hd__nand2_1 _16702_ (.A(_07869_),
    .B(_07870_),
    .Y(_07871_));
 sky130_fd_sc_hd__a21oi_1 _16703_ (.A1(_07778_),
    .A2(_07789_),
    .B1(_07776_),
    .Y(_07872_));
 sky130_fd_sc_hd__or2_1 _16704_ (.A(_07871_),
    .B(_07872_),
    .X(_07873_));
 sky130_fd_sc_hd__nand2_1 _16705_ (.A(_07871_),
    .B(_07872_),
    .Y(_07874_));
 sky130_fd_sc_hd__and2_2 _16706_ (.A(_07873_),
    .B(_07874_),
    .X(_07875_));
 sky130_fd_sc_hd__a21oi_4 _16707_ (.A1(_07695_),
    .A2(_07787_),
    .B1(_07786_),
    .Y(_07876_));
 sky130_fd_sc_hd__nand2b_1 _16708_ (.A_N(_07876_),
    .B(_07875_),
    .Y(_07877_));
 sky130_fd_sc_hd__xnor2_2 _16709_ (.A(_07875_),
    .B(_07876_),
    .Y(_07878_));
 sky130_fd_sc_hd__o21ai_4 _16710_ (.A1(_07791_),
    .A2(_07796_),
    .B1(_07878_),
    .Y(_07880_));
 sky130_fd_sc_hd__or3_1 _16711_ (.A(_07791_),
    .B(_07796_),
    .C(_07878_),
    .X(_07881_));
 sky130_fd_sc_hd__and2_1 _16712_ (.A(_07880_),
    .B(_07881_),
    .X(_07882_));
 sky130_fd_sc_hd__nand2_2 _16713_ (.A(_07798_),
    .B(_07882_),
    .Y(_07883_));
 sky130_fd_sc_hd__or2_1 _16714_ (.A(_07798_),
    .B(_07882_),
    .X(_07884_));
 sky130_fd_sc_hd__nand2_1 _16715_ (.A(_07883_),
    .B(_07884_),
    .Y(_07885_));
 sky130_fd_sc_hd__a21oi_4 _16716_ (.A1(_07712_),
    .A2(_07714_),
    .B1(_07800_),
    .Y(_07886_));
 sky130_fd_sc_hd__a21oi_2 _16717_ (.A1(_07723_),
    .A2(_07801_),
    .B1(_07886_),
    .Y(_07887_));
 sky130_fd_sc_hd__o21ai_1 _16718_ (.A1(_07885_),
    .A2(_07887_),
    .B1(net280),
    .Y(_07888_));
 sky130_fd_sc_hd__a21oi_1 _16719_ (.A1(_07885_),
    .A2(_07887_),
    .B1(_07888_),
    .Y(_07889_));
 sky130_fd_sc_hd__a21bo_1 _16720_ (.A1(net394),
    .A2(net275),
    .B1_N(net701),
    .X(_07891_));
 sky130_fd_sc_hd__inv_2 _16721_ (.A(_07891_),
    .Y(_07892_));
 sky130_fd_sc_hd__nor2_1 _16722_ (.A(net701),
    .B(net271),
    .Y(_07893_));
 sky130_fd_sc_hd__nand2_1 _16723_ (.A(net394),
    .B(_07893_),
    .Y(_07894_));
 sky130_fd_sc_hd__a221o_1 _16724_ (.A1(_07807_),
    .A2(_07810_),
    .B1(_07893_),
    .B2(net394),
    .C1(_07892_),
    .X(_07895_));
 sky130_fd_sc_hd__a211o_1 _16725_ (.A1(_07891_),
    .A2(_07894_),
    .B1(_07806_),
    .C1(_07811_),
    .X(_07896_));
 sky130_fd_sc_hd__a31oi_2 _16726_ (.A1(_02513_),
    .A2(_02551_),
    .A3(_02554_),
    .B1(_02557_),
    .Y(_07897_));
 sky130_fd_sc_hd__nand2b_2 _16727_ (.A_N(_07897_),
    .B(_02543_),
    .Y(_07898_));
 sky130_fd_sc_hd__nand2b_1 _16728_ (.A_N(_02543_),
    .B(_07897_),
    .Y(_07899_));
 sky130_fd_sc_hd__nand2b_1 _16729_ (.A_N(_04334_),
    .B(_05771_),
    .Y(_07900_));
 sky130_fd_sc_hd__xnor2_1 _16730_ (.A(_05822_),
    .B(_07900_),
    .Y(_07902_));
 sky130_fd_sc_hd__a21oi_1 _16731_ (.A1(net697),
    .A2(_05870_),
    .B1(net249),
    .Y(_07903_));
 sky130_fd_sc_hd__o21a_1 _16732_ (.A1(net697),
    .A2(_05870_),
    .B1(_07903_),
    .X(_07904_));
 sky130_fd_sc_hd__a221o_1 _16733_ (.A1(_05771_),
    .A2(net238),
    .B1(net233),
    .B2(net697),
    .C1(net244),
    .X(_07905_));
 sky130_fd_sc_hd__a21o_1 _16734_ (.A1(_04334_),
    .A2(net236),
    .B1(_07905_),
    .X(_07906_));
 sky130_fd_sc_hd__nor2_1 _16735_ (.A(net209),
    .B(_05323_),
    .Y(_07907_));
 sky130_fd_sc_hd__a211o_1 _16736_ (.A1(_05938_),
    .A2(_06359_),
    .B1(_07906_),
    .C1(_07907_),
    .X(_07908_));
 sky130_fd_sc_hd__a211o_4 _16737_ (.A1(net254),
    .A2(_07902_),
    .B1(_07904_),
    .C1(_07908_),
    .X(_07909_));
 sky130_fd_sc_hd__a31o_4 _16738_ (.A1(net260),
    .A2(_07898_),
    .A3(_07899_),
    .B1(_07909_),
    .X(_07910_));
 sky130_fd_sc_hd__a31o_1 _16739_ (.A1(net230),
    .A2(_07895_),
    .A3(_07896_),
    .B1(_07910_),
    .X(_07911_));
 sky130_fd_sc_hd__o2bb2a_2 _16740_ (.A1_N(net701),
    .A2_N(net247),
    .B1(_07889_),
    .B2(_07911_),
    .X(_08698_));
 sky130_fd_sc_hd__o21ai_1 _16741_ (.A1(_07885_),
    .A2(_07887_),
    .B1(_07883_),
    .Y(_07913_));
 sky130_fd_sc_hd__o22a_1 _16742_ (.A1(_06733_),
    .A2(net171),
    .B1(net169),
    .B2(net175),
    .X(_07914_));
 sky130_fd_sc_hd__and4_1 _16743_ (.A(net177),
    .B(net173),
    .C(net172),
    .D(net170),
    .X(_07915_));
 sky130_fd_sc_hd__nor2_2 _16744_ (.A(_07914_),
    .B(_07915_),
    .Y(_07916_));
 sky130_fd_sc_hd__nand2_1 _16745_ (.A(net798),
    .B(net224),
    .Y(_07917_));
 sky130_fd_sc_hd__xnor2_2 _16746_ (.A(_07916_),
    .B(_07917_),
    .Y(_07918_));
 sky130_fd_sc_hd__nor2_4 _16747_ (.A(net183),
    .B(_07009_),
    .Y(_07919_));
 sky130_fd_sc_hd__or3_2 _16748_ (.A(net187),
    .B(net168),
    .C(_07753_),
    .X(_07920_));
 sky130_fd_sc_hd__xnor2_2 _16749_ (.A(_07919_),
    .B(_07920_),
    .Y(_07921_));
 sky130_fd_sc_hd__xnor2_2 _16750_ (.A(_07918_),
    .B(_07921_),
    .Y(_07923_));
 sky130_fd_sc_hd__and3_1 _16751_ (.A(_07836_),
    .B(_07838_),
    .C(_07923_),
    .X(_07924_));
 sky130_fd_sc_hd__a21oi_2 _16752_ (.A1(_07836_),
    .A2(_07838_),
    .B1(_07923_),
    .Y(_07925_));
 sky130_fd_sc_hd__or2_1 _16753_ (.A(_07924_),
    .B(_07925_),
    .X(_07926_));
 sky130_fd_sc_hd__o21a_1 _16754_ (.A1(_07847_),
    .A2(_07850_),
    .B1(_07848_),
    .X(_07927_));
 sky130_fd_sc_hd__o21ai_2 _16755_ (.A1(_07826_),
    .A2(_07829_),
    .B1(_07827_),
    .Y(_07928_));
 sky130_fd_sc_hd__nor2_2 _16756_ (.A(net185),
    .B(_07048_),
    .Y(_07929_));
 sky130_fd_sc_hd__a21oi_1 _16757_ (.A1(net784),
    .A2(net182),
    .B1(_07929_),
    .Y(_07930_));
 sky130_fd_sc_hd__and3_1 _16758_ (.A(net784),
    .B(net182),
    .C(_07929_),
    .X(_07931_));
 sky130_fd_sc_hd__nor2_2 _16759_ (.A(_07930_),
    .B(_07931_),
    .Y(_07932_));
 sky130_fd_sc_hd__nand2_1 _16760_ (.A(net765),
    .B(net132),
    .Y(_07934_));
 sky130_fd_sc_hd__xnor2_2 _16761_ (.A(_07932_),
    .B(_07934_),
    .Y(_07935_));
 sky130_fd_sc_hd__xor2_1 _16762_ (.A(_07928_),
    .B(_07935_),
    .X(_07936_));
 sky130_fd_sc_hd__and2b_1 _16763_ (.A_N(_07927_),
    .B(_07936_),
    .X(_07937_));
 sky130_fd_sc_hd__and2b_1 _16764_ (.A_N(_07936_),
    .B(_07927_),
    .X(_07938_));
 sky130_fd_sc_hd__or2_1 _16765_ (.A(_07937_),
    .B(_07938_),
    .X(_07939_));
 sky130_fd_sc_hd__and2_1 _16766_ (.A(_07926_),
    .B(_07939_),
    .X(_07940_));
 sky130_fd_sc_hd__nor2_1 _16767_ (.A(_07926_),
    .B(_07939_),
    .Y(_07941_));
 sky130_fd_sc_hd__nor2_1 _16768_ (.A(_07940_),
    .B(_07941_),
    .Y(_07942_));
 sky130_fd_sc_hd__o21ai_1 _16769_ (.A1(_07842_),
    .A2(_07856_),
    .B1(_07942_),
    .Y(_07943_));
 sky130_fd_sc_hd__or3_1 _16770_ (.A(_07842_),
    .B(_07856_),
    .C(_07942_),
    .X(_07945_));
 sky130_fd_sc_hd__and2_2 _16771_ (.A(_07943_),
    .B(_07945_),
    .X(_07946_));
 sky130_fd_sc_hd__a21o_1 _16772_ (.A1(_07845_),
    .A2(_07853_),
    .B1(_07852_),
    .X(_07947_));
 sky130_fd_sc_hd__and2b_1 _16773_ (.A_N(_07780_),
    .B(_07947_),
    .X(_07948_));
 sky130_fd_sc_hd__xnor2_2 _16774_ (.A(_07780_),
    .B(_07947_),
    .Y(_07949_));
 sky130_fd_sc_hd__xnor2_2 _16775_ (.A(_07946_),
    .B(_07949_),
    .Y(_07950_));
 sky130_fd_sc_hd__a21oi_2 _16776_ (.A1(_07860_),
    .A2(_07869_),
    .B1(_07950_),
    .Y(_07951_));
 sky130_fd_sc_hd__and3_1 _16777_ (.A(_07860_),
    .B(_07869_),
    .C(_07950_),
    .X(_07952_));
 sky130_fd_sc_hd__or2_1 _16778_ (.A(_07951_),
    .B(_07952_),
    .X(_07953_));
 sky130_fd_sc_hd__a21boi_1 _16779_ (.A1(_07783_),
    .A2(_07865_),
    .B1_N(_07864_),
    .Y(_07954_));
 sky130_fd_sc_hd__nor2_1 _16780_ (.A(_07953_),
    .B(_07954_),
    .Y(_07956_));
 sky130_fd_sc_hd__and2_1 _16781_ (.A(_07953_),
    .B(_07954_),
    .X(_07957_));
 sky130_fd_sc_hd__or2_1 _16782_ (.A(_07956_),
    .B(_07957_),
    .X(_07958_));
 sky130_fd_sc_hd__a21oi_2 _16783_ (.A1(_07873_),
    .A2(_07877_),
    .B1(_07958_),
    .Y(_07959_));
 sky130_fd_sc_hd__and3_1 _16784_ (.A(_07873_),
    .B(_07877_),
    .C(_07958_),
    .X(_07960_));
 sky130_fd_sc_hd__or2_2 _16785_ (.A(_07959_),
    .B(_07960_),
    .X(_07961_));
 sky130_fd_sc_hd__xor2_2 _16786_ (.A(_07880_),
    .B(_07961_),
    .X(_07962_));
 sky130_fd_sc_hd__xnor2_1 _16787_ (.A(_07913_),
    .B(_07962_),
    .Y(_07963_));
 sky130_fd_sc_hd__a21boi_2 _16788_ (.A1(net385),
    .A2(net274),
    .B1_N(net691),
    .Y(_07964_));
 sky130_fd_sc_hd__nor2_1 _16789_ (.A(net691),
    .B(net271),
    .Y(_07965_));
 sky130_fd_sc_hd__a21oi_2 _16790_ (.A1(net385),
    .A2(_07965_),
    .B1(_07964_),
    .Y(_07967_));
 sky130_fd_sc_hd__nand2_1 _16791_ (.A(_07891_),
    .B(_07895_),
    .Y(_07968_));
 sky130_fd_sc_hd__xnor2_1 _16792_ (.A(_07967_),
    .B(_07968_),
    .Y(_07969_));
 sky130_fd_sc_hd__or2_1 _16793_ (.A(net229),
    .B(_07969_),
    .X(_07970_));
 sky130_fd_sc_hd__nand2_2 _16794_ (.A(_02541_),
    .B(_07898_),
    .Y(_07971_));
 sky130_fd_sc_hd__xnor2_4 _16795_ (.A(_02545_),
    .B(_07971_),
    .Y(_07972_));
 sky130_fd_sc_hd__nand2_1 _16796_ (.A(_04597_),
    .B(_05770_),
    .Y(_07973_));
 sky130_fd_sc_hd__xor2_1 _16797_ (.A(_05824_),
    .B(_07973_),
    .X(_07974_));
 sky130_fd_sc_hd__a21oi_1 _16798_ (.A1(net697),
    .A2(_05870_),
    .B1(net688),
    .Y(_07975_));
 sky130_fd_sc_hd__a221o_1 _16799_ (.A1(_05770_),
    .A2(net238),
    .B1(net233),
    .B2(net688),
    .C1(net244),
    .X(_07976_));
 sky130_fd_sc_hd__a31o_1 _16800_ (.A1(net386),
    .A2(net688),
    .A3(net236),
    .B1(_07976_),
    .X(_07978_));
 sky130_fd_sc_hd__a21oi_1 _16801_ (.A1(_05938_),
    .A2(_06437_),
    .B1(_07978_),
    .Y(_07979_));
 sky130_fd_sc_hd__o21a_1 _16802_ (.A1(net211),
    .A2(_05394_),
    .B1(_07979_),
    .X(_07980_));
 sky130_fd_sc_hd__o31a_1 _16803_ (.A1(net249),
    .A2(_05871_),
    .A3(_07975_),
    .B1(_07980_),
    .X(_07981_));
 sky130_fd_sc_hd__o221a_2 _16804_ (.A1(net257),
    .A2(_07972_),
    .B1(_07974_),
    .B2(net253),
    .C1(_07981_),
    .X(_07982_));
 sky130_fd_sc_hd__o211a_1 _16805_ (.A1(net278),
    .A2(_07963_),
    .B1(_07970_),
    .C1(_07982_),
    .X(_07983_));
 sky130_fd_sc_hd__a21oi_2 _16806_ (.A1(net691),
    .A2(net246),
    .B1(_07983_),
    .Y(_08699_));
 sky130_fd_sc_hd__nand2_1 _16807_ (.A(net784),
    .B(net223),
    .Y(_07984_));
 sky130_fd_sc_hd__a22o_1 _16808_ (.A1(net472),
    .A2(net173),
    .B1(net172),
    .B2(net797),
    .X(_07985_));
 sky130_fd_sc_hd__and3_1 _16809_ (.A(net472),
    .B(_00653_),
    .C(net173),
    .X(_07986_));
 sky130_fd_sc_hd__o31a_1 _16810_ (.A1(_00654_),
    .A2(_06733_),
    .A3(net169),
    .B1(_07985_),
    .X(_07988_));
 sky130_fd_sc_hd__xnor2_1 _16811_ (.A(_07984_),
    .B(_07988_),
    .Y(_07989_));
 sky130_fd_sc_hd__or4b_1 _16812_ (.A(net188),
    .B(net175),
    .C(net168),
    .D_N(_07919_),
    .X(_07990_));
 sky130_fd_sc_hd__nor2_1 _16813_ (.A(net175),
    .B(_07009_),
    .Y(_07991_));
 sky130_fd_sc_hd__or4b_2 _16814_ (.A(net187),
    .B(net177),
    .C(net168),
    .D_N(_07919_),
    .X(_07992_));
 sky130_fd_sc_hd__a21o_1 _16815_ (.A1(net452),
    .A2(net184),
    .B1(_07991_),
    .X(_07993_));
 sky130_fd_sc_hd__and3_1 _16816_ (.A(_07990_),
    .B(_07992_),
    .C(_07993_),
    .X(_07994_));
 sky130_fd_sc_hd__or2_1 _16817_ (.A(_07989_),
    .B(_07994_),
    .X(_07995_));
 sky130_fd_sc_hd__nand2_1 _16818_ (.A(_07989_),
    .B(_07994_),
    .Y(_07996_));
 sky130_fd_sc_hd__nand2_1 _16819_ (.A(_07995_),
    .B(_07996_),
    .Y(_07997_));
 sky130_fd_sc_hd__o2bb2a_1 _16820_ (.A1_N(_07918_),
    .A2_N(_07921_),
    .B1(_07919_),
    .B2(_07832_),
    .X(_07999_));
 sky130_fd_sc_hd__nor2_1 _16821_ (.A(_07997_),
    .B(_07999_),
    .Y(_08000_));
 sky130_fd_sc_hd__and2_1 _16822_ (.A(_07997_),
    .B(_07999_),
    .X(_08001_));
 sky130_fd_sc_hd__or2_1 _16823_ (.A(_08000_),
    .B(_08001_),
    .X(_08002_));
 sky130_fd_sc_hd__a31o_1 _16824_ (.A1(net765),
    .A2(net132),
    .A3(_07932_),
    .B1(_07931_),
    .X(_08003_));
 sky130_fd_sc_hd__a31o_2 _16825_ (.A1(net797),
    .A2(net224),
    .A3(_07916_),
    .B1(_07915_),
    .X(_08004_));
 sky130_fd_sc_hd__a22o_1 _16826_ (.A1(net776),
    .A2(net182),
    .B1(_07164_),
    .B2(_06530_),
    .X(_08005_));
 sky130_fd_sc_hd__or4_2 _16827_ (.A(net185),
    .B(net179),
    .C(_07048_),
    .D(_07165_),
    .X(_08006_));
 sky130_fd_sc_hd__nand2_1 _16828_ (.A(_08005_),
    .B(_08006_),
    .Y(_08007_));
 sky130_fd_sc_hd__xnor2_2 _16829_ (.A(_08004_),
    .B(_08007_),
    .Y(_08008_));
 sky130_fd_sc_hd__xnor2_1 _16830_ (.A(_08003_),
    .B(_08008_),
    .Y(_08010_));
 sky130_fd_sc_hd__and2_1 _16831_ (.A(_08002_),
    .B(_08010_),
    .X(_08011_));
 sky130_fd_sc_hd__nor2_1 _16832_ (.A(_08002_),
    .B(_08010_),
    .Y(_08012_));
 sky130_fd_sc_hd__nor2_1 _16833_ (.A(_08011_),
    .B(_08012_),
    .Y(_08013_));
 sky130_fd_sc_hd__o21a_1 _16834_ (.A1(_07925_),
    .A2(_07941_),
    .B1(_08013_),
    .X(_08014_));
 sky130_fd_sc_hd__nor3_1 _16835_ (.A(_07925_),
    .B(_07941_),
    .C(_08013_),
    .Y(_08015_));
 sky130_fd_sc_hd__nor2_2 _16836_ (.A(_08014_),
    .B(_08015_),
    .Y(_08016_));
 sky130_fd_sc_hd__a21o_1 _16837_ (.A1(_07928_),
    .A2(_07935_),
    .B1(_07937_),
    .X(_08017_));
 sky130_fd_sc_hd__xnor2_2 _16838_ (.A(_08016_),
    .B(_08017_),
    .Y(_08018_));
 sky130_fd_sc_hd__a21bo_1 _16839_ (.A1(_07946_),
    .A2(_07949_),
    .B1_N(_07943_),
    .X(_08019_));
 sky130_fd_sc_hd__nand2b_1 _16840_ (.A_N(_08018_),
    .B(_08019_),
    .Y(_08021_));
 sky130_fd_sc_hd__xnor2_1 _16841_ (.A(_08018_),
    .B(_08019_),
    .Y(_08022_));
 sky130_fd_sc_hd__nand2_1 _16842_ (.A(_07948_),
    .B(_08022_),
    .Y(_08023_));
 sky130_fd_sc_hd__or2_1 _16843_ (.A(_07948_),
    .B(_08022_),
    .X(_08024_));
 sky130_fd_sc_hd__and2_1 _16844_ (.A(_08023_),
    .B(_08024_),
    .X(_08025_));
 sky130_fd_sc_hd__o21ai_2 _16845_ (.A1(_07951_),
    .A2(_07956_),
    .B1(_08025_),
    .Y(_08026_));
 sky130_fd_sc_hd__or3_1 _16846_ (.A(_07951_),
    .B(_07956_),
    .C(_08025_),
    .X(_08027_));
 sky130_fd_sc_hd__nand2_1 _16847_ (.A(_08026_),
    .B(_08027_),
    .Y(_08028_));
 sky130_fd_sc_hd__inv_2 _16848_ (.A(_08028_),
    .Y(_08029_));
 sky130_fd_sc_hd__nand2_1 _16849_ (.A(_07959_),
    .B(_08029_),
    .Y(_08030_));
 sky130_fd_sc_hd__or2_1 _16850_ (.A(_07959_),
    .B(_08029_),
    .X(_08032_));
 sky130_fd_sc_hd__nand2_1 _16851_ (.A(_08030_),
    .B(_08032_),
    .Y(_08033_));
 sky130_fd_sc_hd__a21oi_2 _16852_ (.A1(_07880_),
    .A2(_07883_),
    .B1(_07961_),
    .Y(_08034_));
 sky130_fd_sc_hd__and3_2 _16853_ (.A(_07883_),
    .B(_07884_),
    .C(_07962_),
    .X(_08035_));
 sky130_fd_sc_hd__and4bb_2 _16854_ (.A_N(_07717_),
    .B_N(_07722_),
    .C(_07801_),
    .D(_08035_),
    .X(_08036_));
 sky130_fd_sc_hd__a211oi_4 _16855_ (.A1(_07886_),
    .A2(_08035_),
    .B1(_08036_),
    .C1(_08034_),
    .Y(_08037_));
 sky130_fd_sc_hd__o21ai_1 _16856_ (.A1(_08033_),
    .A2(_08037_),
    .B1(net280),
    .Y(_08038_));
 sky130_fd_sc_hd__a21oi_1 _16857_ (.A1(_08033_),
    .A2(_08037_),
    .B1(_08038_),
    .Y(_08039_));
 sky130_fd_sc_hd__a21boi_4 _16858_ (.A1(net378),
    .A2(net274),
    .B1_N(net681),
    .Y(_08040_));
 sky130_fd_sc_hd__nor2_1 _16859_ (.A(net681),
    .B(_05955_),
    .Y(_08041_));
 sky130_fd_sc_hd__a21oi_4 _16860_ (.A1(net378),
    .A2(_08041_),
    .B1(_08040_),
    .Y(_08043_));
 sky130_fd_sc_hd__a21o_2 _16861_ (.A1(_07967_),
    .A2(_07968_),
    .B1(_07964_),
    .X(_08044_));
 sky130_fd_sc_hd__or2_1 _16862_ (.A(_08043_),
    .B(_08044_),
    .X(_08045_));
 sky130_fd_sc_hd__nand2_1 _16863_ (.A(_08043_),
    .B(_08044_),
    .Y(_08046_));
 sky130_fd_sc_hd__nand2_1 _16864_ (.A(_04820_),
    .B(_05769_),
    .Y(_08047_));
 sky130_fd_sc_hd__xnor2_1 _16865_ (.A(_05825_),
    .B(_08047_),
    .Y(_08048_));
 sky130_fd_sc_hd__nand2_1 _16866_ (.A(_01579_),
    .B(_02560_),
    .Y(_08049_));
 sky130_fd_sc_hd__o21ai_1 _16867_ (.A1(net678),
    .A2(_05871_),
    .B1(_05849_),
    .Y(_08050_));
 sky130_fd_sc_hd__nor2_1 _16868_ (.A(_05872_),
    .B(_08050_),
    .Y(_08051_));
 sky130_fd_sc_hd__a221o_1 _16869_ (.A1(_05769_),
    .A2(net238),
    .B1(net233),
    .B2(net678),
    .C1(net244),
    .X(_08052_));
 sky130_fd_sc_hd__a31o_1 _16870_ (.A1(net379),
    .A2(net679),
    .A3(net236),
    .B1(_08052_),
    .X(_08054_));
 sky130_fd_sc_hd__o22a_1 _16871_ (.A1(net210),
    .A2(_05459_),
    .B1(net203),
    .B2(_06519_),
    .X(_08055_));
 sky130_fd_sc_hd__or3b_4 _16872_ (.A(_08051_),
    .B(_08054_),
    .C_N(_08055_),
    .X(_08056_));
 sky130_fd_sc_hd__a31o_2 _16873_ (.A1(_02561_),
    .A2(net260),
    .A3(_08049_),
    .B1(_08056_),
    .X(_08057_));
 sky130_fd_sc_hd__a21o_2 _16874_ (.A1(_05840_),
    .A2(_08048_),
    .B1(_08057_),
    .X(_08058_));
 sky130_fd_sc_hd__a31o_1 _16875_ (.A1(net230),
    .A2(_08045_),
    .A3(_08046_),
    .B1(_08058_),
    .X(_08059_));
 sky130_fd_sc_hd__o2bb2a_2 _16876_ (.A1_N(net681),
    .A2_N(net246),
    .B1(_08039_),
    .B2(_08059_),
    .X(_08700_));
 sky130_fd_sc_hd__o21ai_1 _16877_ (.A1(_08033_),
    .A2(_08037_),
    .B1(_08030_),
    .Y(_08060_));
 sky130_fd_sc_hd__a21o_1 _16878_ (.A1(net468),
    .A2(net793),
    .B1(_00506_),
    .X(_08061_));
 sky130_fd_sc_hd__o211a_4 _16879_ (.A1(_00220_),
    .A2(_00654_),
    .B1(_06179_),
    .C1(_08061_),
    .X(_08062_));
 sky130_fd_sc_hd__and3_2 _16880_ (.A(net775),
    .B(net223),
    .C(_08062_),
    .X(_08064_));
 sky130_fd_sc_hd__a21oi_1 _16881_ (.A1(net775),
    .A2(net223),
    .B1(_08062_),
    .Y(_08065_));
 sky130_fd_sc_hd__or2_1 _16882_ (.A(_08064_),
    .B(_08065_),
    .X(_08066_));
 sky130_fd_sc_hd__or3_1 _16883_ (.A(net175),
    .B(net168),
    .C(_07919_),
    .X(_08067_));
 sky130_fd_sc_hd__xnor2_1 _16884_ (.A(_07010_),
    .B(_08067_),
    .Y(_08068_));
 sky130_fd_sc_hd__nor2_1 _16885_ (.A(_08066_),
    .B(_08068_),
    .Y(_08069_));
 sky130_fd_sc_hd__and2_1 _16886_ (.A(_08066_),
    .B(_08068_),
    .X(_08070_));
 sky130_fd_sc_hd__or2_1 _16887_ (.A(_08069_),
    .B(_08070_),
    .X(_08071_));
 sky130_fd_sc_hd__nand3_1 _16888_ (.A(_07992_),
    .B(_07996_),
    .C(_08071_),
    .Y(_08072_));
 sky130_fd_sc_hd__a21o_2 _16889_ (.A1(_07992_),
    .A2(_07996_),
    .B1(_08071_),
    .X(_08073_));
 sky130_fd_sc_hd__nand2_1 _16890_ (.A(_08072_),
    .B(_08073_),
    .Y(_08075_));
 sky130_fd_sc_hd__a31o_1 _16891_ (.A1(net784),
    .A2(net223),
    .A3(_07985_),
    .B1(_07986_),
    .X(_08076_));
 sky130_fd_sc_hd__o211a_1 _16892_ (.A1(net185),
    .A2(_07048_),
    .B1(net182),
    .C1(net762),
    .X(_08077_));
 sky130_fd_sc_hd__xnor2_1 _16893_ (.A(_08076_),
    .B(_08077_),
    .Y(_08078_));
 sky130_fd_sc_hd__or2_2 _16894_ (.A(_08075_),
    .B(_08078_),
    .X(_08079_));
 sky130_fd_sc_hd__nand2_1 _16895_ (.A(_08075_),
    .B(_08078_),
    .Y(_08080_));
 sky130_fd_sc_hd__and2_1 _16896_ (.A(_08079_),
    .B(_08080_),
    .X(_08081_));
 sky130_fd_sc_hd__or3_2 _16897_ (.A(_08000_),
    .B(_08012_),
    .C(_08081_),
    .X(_08082_));
 sky130_fd_sc_hd__o21ai_2 _16898_ (.A1(_08000_),
    .A2(_08012_),
    .B1(_08081_),
    .Y(_08083_));
 sky130_fd_sc_hd__a32o_2 _16899_ (.A1(_08004_),
    .A2(_08005_),
    .A3(_08006_),
    .B1(_08008_),
    .B2(_08003_),
    .X(_08084_));
 sky130_fd_sc_hd__and3_1 _16900_ (.A(_08082_),
    .B(_08083_),
    .C(_08084_),
    .X(_08086_));
 sky130_fd_sc_hd__a21oi_2 _16901_ (.A1(_08082_),
    .A2(_08083_),
    .B1(_08084_),
    .Y(_08087_));
 sky130_fd_sc_hd__nor2_4 _16902_ (.A(_08086_),
    .B(_08087_),
    .Y(_08088_));
 sky130_fd_sc_hd__a21o_2 _16903_ (.A1(_08016_),
    .A2(_08017_),
    .B1(_08014_),
    .X(_08089_));
 sky130_fd_sc_hd__nand2_1 _16904_ (.A(_08088_),
    .B(_08089_),
    .Y(_08090_));
 sky130_fd_sc_hd__xnor2_4 _16905_ (.A(_08088_),
    .B(_08089_),
    .Y(_08091_));
 sky130_fd_sc_hd__nand2_1 _16906_ (.A(_08021_),
    .B(_08023_),
    .Y(_08092_));
 sky130_fd_sc_hd__a21o_1 _16907_ (.A1(_08021_),
    .A2(_08023_),
    .B1(_08091_),
    .X(_08093_));
 sky130_fd_sc_hd__xnor2_2 _16908_ (.A(_08091_),
    .B(_08092_),
    .Y(_08094_));
 sky130_fd_sc_hd__xnor2_1 _16909_ (.A(_08026_),
    .B(_08094_),
    .Y(_08095_));
 sky130_fd_sc_hd__xor2_1 _16910_ (.A(_08060_),
    .B(_08095_),
    .X(_08097_));
 sky130_fd_sc_hd__nand2_2 _16911_ (.A(net280),
    .B(_08097_),
    .Y(_08098_));
 sky130_fd_sc_hd__a21boi_2 _16912_ (.A1(net369),
    .A2(net275),
    .B1_N(net672),
    .Y(_08099_));
 sky130_fd_sc_hd__and3b_1 _16913_ (.A_N(net672),
    .B(net274),
    .C(net369),
    .X(_08100_));
 sky130_fd_sc_hd__nor2_2 _16914_ (.A(_08099_),
    .B(_08100_),
    .Y(_08101_));
 sky130_fd_sc_hd__a21oi_1 _16915_ (.A1(_08043_),
    .A2(_08044_),
    .B1(_08040_),
    .Y(_08102_));
 sky130_fd_sc_hd__xnor2_1 _16916_ (.A(_08101_),
    .B(_08102_),
    .Y(_08103_));
 sky130_fd_sc_hd__nand2_1 _16917_ (.A(net230),
    .B(_08103_),
    .Y(_08104_));
 sky130_fd_sc_hd__and3_1 _16918_ (.A(_04929_),
    .B(_05767_),
    .C(_05826_),
    .X(_08105_));
 sky130_fd_sc_hd__a21oi_1 _16919_ (.A1(_04929_),
    .A2(_05767_),
    .B1(_05826_),
    .Y(_08106_));
 sky130_fd_sc_hd__o21ai_1 _16920_ (.A1(_01483_),
    .A2(_01576_),
    .B1(_02561_),
    .Y(_08108_));
 sky130_fd_sc_hd__xnor2_1 _16921_ (.A(_02563_),
    .B(_08108_),
    .Y(_08109_));
 sky130_fd_sc_hd__nand2_2 _16922_ (.A(net260),
    .B(_08109_),
    .Y(_08110_));
 sky130_fd_sc_hd__a21oi_1 _16923_ (.A1(net674),
    .A2(_05872_),
    .B1(net250),
    .Y(_08111_));
 sky130_fd_sc_hd__o21ai_1 _16924_ (.A1(net674),
    .A2(_05872_),
    .B1(_08111_),
    .Y(_08112_));
 sky130_fd_sc_hd__a221o_1 _16925_ (.A1(_05767_),
    .A2(net238),
    .B1(net233),
    .B2(net674),
    .C1(net244),
    .X(_08113_));
 sky130_fd_sc_hd__a21oi_1 _16926_ (.A1(_04928_),
    .A2(net236),
    .B1(_08113_),
    .Y(_08114_));
 sky130_fd_sc_hd__o21a_1 _16927_ (.A1(_05939_),
    .A2(_06602_),
    .B1(_08114_),
    .X(_08115_));
 sky130_fd_sc_hd__o211a_1 _16928_ (.A1(net548),
    .A2(_05525_),
    .B1(_08112_),
    .C1(_08115_),
    .X(_08116_));
 sky130_fd_sc_hd__o311a_4 _16929_ (.A1(net252),
    .A2(_08105_),
    .A3(_08106_),
    .B1(_08110_),
    .C1(_08116_),
    .X(_08117_));
 sky130_fd_sc_hd__a32oi_4 _16930_ (.A1(_08098_),
    .A2(_08104_),
    .A3(_08117_),
    .B1(net246),
    .B2(net672),
    .Y(_08701_));
 sky130_fd_sc_hd__or3b_2 _16931_ (.A(_08033_),
    .B(_08037_),
    .C_N(_08095_),
    .X(_08119_));
 sky130_fd_sc_hd__a21bo_1 _16932_ (.A1(_08026_),
    .A2(_08030_),
    .B1_N(_08094_),
    .X(_08120_));
 sky130_fd_sc_hd__nand2_1 _16933_ (.A(_00220_),
    .B(_00363_),
    .Y(_08121_));
 sky130_fd_sc_hd__o211a_4 _16934_ (.A1(_08625_),
    .A2(_00507_),
    .B1(_06179_),
    .C1(_08121_),
    .X(_08122_));
 sky130_fd_sc_hd__and3_1 _16935_ (.A(net762),
    .B(net223),
    .C(_08122_),
    .X(_08123_));
 sky130_fd_sc_hd__a21oi_1 _16936_ (.A1(net762),
    .A2(net223),
    .B1(_08122_),
    .Y(_08124_));
 sky130_fd_sc_hd__nor2_1 _16937_ (.A(_08123_),
    .B(_08124_),
    .Y(_08125_));
 sky130_fd_sc_hd__or4_1 _16938_ (.A(net797),
    .B(net175),
    .C(_07010_),
    .D(net168),
    .X(_08126_));
 sky130_fd_sc_hd__or2_2 _16939_ (.A(_00207_),
    .B(_07010_),
    .X(_08127_));
 sky130_fd_sc_hd__a22o_1 _16940_ (.A1(net461),
    .A2(_06827_),
    .B1(_07128_),
    .B2(net173),
    .X(_08129_));
 sky130_fd_sc_hd__o211a_1 _16941_ (.A1(_07991_),
    .A2(_08127_),
    .B1(_08129_),
    .C1(_08126_),
    .X(_08130_));
 sky130_fd_sc_hd__nand2_1 _16942_ (.A(_08125_),
    .B(_08130_),
    .Y(_08131_));
 sky130_fd_sc_hd__or2_2 _16943_ (.A(_08125_),
    .B(_08130_),
    .X(_08132_));
 sky130_fd_sc_hd__nand2_4 _16944_ (.A(_08131_),
    .B(_08132_),
    .Y(_08133_));
 sky130_fd_sc_hd__a41o_4 _16945_ (.A1(net177),
    .A2(_06733_),
    .A3(_07128_),
    .A4(_07919_),
    .B1(_08069_),
    .X(_08134_));
 sky130_fd_sc_hd__nand2b_1 _16946_ (.A_N(_08133_),
    .B(_08134_),
    .Y(_08135_));
 sky130_fd_sc_hd__xnor2_4 _16947_ (.A(_08133_),
    .B(_08134_),
    .Y(_08136_));
 sky130_fd_sc_hd__a31oi_4 _16948_ (.A1(net797),
    .A2(_00219_),
    .A3(net172),
    .B1(_08064_),
    .Y(_08137_));
 sky130_fd_sc_hd__nand2b_1 _16949_ (.A_N(_08137_),
    .B(_08136_),
    .Y(_08138_));
 sky130_fd_sc_hd__xor2_4 _16950_ (.A(_08136_),
    .B(_08137_),
    .X(_08140_));
 sky130_fd_sc_hd__a21oi_4 _16951_ (.A1(_08073_),
    .A2(_08079_),
    .B1(_08140_),
    .Y(_08141_));
 sky130_fd_sc_hd__and3_1 _16952_ (.A(_08073_),
    .B(_08079_),
    .C(_08140_),
    .X(_08142_));
 sky130_fd_sc_hd__nor2_4 _16953_ (.A(_08141_),
    .B(_08142_),
    .Y(_08143_));
 sky130_fd_sc_hd__o211a_4 _16954_ (.A1(_07929_),
    .A2(_08076_),
    .B1(net762),
    .C1(net182),
    .X(_08144_));
 sky130_fd_sc_hd__xnor2_4 _16955_ (.A(_08143_),
    .B(_08144_),
    .Y(_08145_));
 sky130_fd_sc_hd__a21bo_2 _16956_ (.A1(_08082_),
    .A2(_08084_),
    .B1_N(_08083_),
    .X(_08146_));
 sky130_fd_sc_hd__nand2b_1 _16957_ (.A_N(_08145_),
    .B(_08146_),
    .Y(_08147_));
 sky130_fd_sc_hd__xor2_4 _16958_ (.A(_08145_),
    .B(_08146_),
    .X(_08148_));
 sky130_fd_sc_hd__nand2_1 _16959_ (.A(_08090_),
    .B(_08093_),
    .Y(_08149_));
 sky130_fd_sc_hd__xor2_1 _16960_ (.A(_08148_),
    .B(_08149_),
    .X(_08151_));
 sky130_fd_sc_hd__a21o_1 _16961_ (.A1(_08119_),
    .A2(_08120_),
    .B1(_08151_),
    .X(_08152_));
 sky130_fd_sc_hd__nand2_1 _16962_ (.A(net281),
    .B(_08152_),
    .Y(_08153_));
 sky130_fd_sc_hd__a31o_1 _16963_ (.A1(_08119_),
    .A2(_08120_),
    .A3(_08151_),
    .B1(_08153_),
    .X(_08154_));
 sky130_fd_sc_hd__a21boi_1 _16964_ (.A1(net360),
    .A2(net274),
    .B1_N(net664),
    .Y(_08155_));
 sky130_fd_sc_hd__and3b_1 _16965_ (.A_N(net664),
    .B(net274),
    .C(net360),
    .X(_08156_));
 sky130_fd_sc_hd__or2_1 _16966_ (.A(_08155_),
    .B(_08156_),
    .X(_08157_));
 sky130_fd_sc_hd__o21ba_1 _16967_ (.A1(_08040_),
    .A2(_08099_),
    .B1_N(_08100_),
    .X(_08158_));
 sky130_fd_sc_hd__a31oi_4 _16968_ (.A1(_08043_),
    .A2(_08044_),
    .A3(_08101_),
    .B1(_08158_),
    .Y(_08159_));
 sky130_fd_sc_hd__xnor2_1 _16969_ (.A(_08157_),
    .B(_08159_),
    .Y(_08160_));
 sky130_fd_sc_hd__nand2_1 _16970_ (.A(_05182_),
    .B(_05766_),
    .Y(_08162_));
 sky130_fd_sc_hd__xnor2_1 _16971_ (.A(_05827_),
    .B(_08162_),
    .Y(_08163_));
 sky130_fd_sc_hd__xnor2_4 _16972_ (.A(_01378_),
    .B(_02564_),
    .Y(_08164_));
 sky130_fd_sc_hd__a21oi_1 _16973_ (.A1(net674),
    .A2(_05872_),
    .B1(net666),
    .Y(_08165_));
 sky130_fd_sc_hd__nand2_1 _16974_ (.A(net666),
    .B(net232),
    .Y(_08166_));
 sky130_fd_sc_hd__o221a_1 _16975_ (.A1(_05765_),
    .A2(_05942_),
    .B1(net235),
    .B2(_05182_),
    .C1(_08166_),
    .X(_08167_));
 sky130_fd_sc_hd__o22a_1 _16976_ (.A1(net211),
    .A2(_05575_),
    .B1(net203),
    .B2(_06700_),
    .X(_08168_));
 sky130_fd_sc_hd__and3_1 _16977_ (.A(_05880_),
    .B(_08167_),
    .C(_08168_),
    .X(_08169_));
 sky130_fd_sc_hd__o31a_1 _16978_ (.A1(net250),
    .A2(_05873_),
    .A3(_08165_),
    .B1(_08169_),
    .X(_08170_));
 sky130_fd_sc_hd__o221a_1 _16979_ (.A1(net252),
    .A2(_08163_),
    .B1(_08164_),
    .B2(net257),
    .C1(_08170_),
    .X(_08171_));
 sky130_fd_sc_hd__o211a_1 _16980_ (.A1(net229),
    .A2(_08160_),
    .B1(_08171_),
    .C1(_08154_),
    .X(_08173_));
 sky130_fd_sc_hd__a21oi_1 _16981_ (.A1(net664),
    .A2(net246),
    .B1(_08173_),
    .Y(_08702_));
 sky130_fd_sc_hd__or3_2 _16982_ (.A(_08613_),
    .B(_00361_),
    .C(net266),
    .X(_08174_));
 sky130_fd_sc_hd__nand2_1 _16983_ (.A(_00207_),
    .B(_00221_),
    .Y(_08175_));
 sky130_fd_sc_hd__and3_1 _16984_ (.A(net227),
    .B(_08174_),
    .C(_08175_),
    .X(_08176_));
 sky130_fd_sc_hd__and2b_1 _16985_ (.A_N(_08127_),
    .B(_08176_),
    .X(_08177_));
 sky130_fd_sc_hd__xnor2_1 _16986_ (.A(_08127_),
    .B(_08176_),
    .Y(_08178_));
 sky130_fd_sc_hd__nand2_1 _16987_ (.A(net762),
    .B(net170),
    .Y(_08179_));
 sky130_fd_sc_hd__nor2_1 _16988_ (.A(_00363_),
    .B(_08179_),
    .Y(_08180_));
 sky130_fd_sc_hd__or2_1 _16989_ (.A(_00363_),
    .B(_08179_),
    .X(_08181_));
 sky130_fd_sc_hd__nand2_4 _16990_ (.A(_08625_),
    .B(_00223_),
    .Y(_08183_));
 sky130_fd_sc_hd__and4_1 _16991_ (.A(net227),
    .B(_08178_),
    .C(_08181_),
    .D(_08183_),
    .X(_08184_));
 sky130_fd_sc_hd__a31o_1 _16992_ (.A1(net227),
    .A2(_08181_),
    .A3(_08183_),
    .B1(_08178_),
    .X(_08185_));
 sky130_fd_sc_hd__and2b_1 _16993_ (.A_N(_08184_),
    .B(_08185_),
    .X(_08186_));
 sky130_fd_sc_hd__and2_1 _16994_ (.A(_08126_),
    .B(_08131_),
    .X(_08187_));
 sky130_fd_sc_hd__and2b_1 _16995_ (.A_N(_08186_),
    .B(_08187_),
    .X(_08188_));
 sky130_fd_sc_hd__and2b_1 _16996_ (.A_N(_08187_),
    .B(_08186_),
    .X(_08189_));
 sky130_fd_sc_hd__nor2_1 _16997_ (.A(_08188_),
    .B(_08189_),
    .Y(_08190_));
 sky130_fd_sc_hd__a31o_1 _16998_ (.A1(net775),
    .A2(_00219_),
    .A3(net172),
    .B1(_08123_),
    .X(_08191_));
 sky130_fd_sc_hd__and2_1 _16999_ (.A(_08190_),
    .B(_08191_),
    .X(_08192_));
 sky130_fd_sc_hd__nor2_1 _17000_ (.A(_08190_),
    .B(_08191_),
    .Y(_08194_));
 sky130_fd_sc_hd__or2_1 _17001_ (.A(_08192_),
    .B(_08194_),
    .X(_08195_));
 sky130_fd_sc_hd__a21o_2 _17002_ (.A1(_08135_),
    .A2(_08138_),
    .B1(_08195_),
    .X(_08196_));
 sky130_fd_sc_hd__nand3_2 _17003_ (.A(_08135_),
    .B(_08138_),
    .C(_08195_),
    .Y(_08197_));
 sky130_fd_sc_hd__nand2_4 _17004_ (.A(_08196_),
    .B(_08197_),
    .Y(_08198_));
 sky130_fd_sc_hd__a21oi_4 _17005_ (.A1(_08143_),
    .A2(_08144_),
    .B1(_08141_),
    .Y(_08199_));
 sky130_fd_sc_hd__or2_1 _17006_ (.A(_08198_),
    .B(_08199_),
    .X(_08200_));
 sky130_fd_sc_hd__xnor2_4 _17007_ (.A(_08198_),
    .B(_08199_),
    .Y(_08201_));
 sky130_fd_sc_hd__or2_2 _17008_ (.A(_08090_),
    .B(_08148_),
    .X(_08202_));
 sky130_fd_sc_hd__nand2_2 _17009_ (.A(_08147_),
    .B(_08202_),
    .Y(_08203_));
 sky130_fd_sc_hd__xor2_4 _17010_ (.A(_08201_),
    .B(_08203_),
    .X(_08205_));
 sky130_fd_sc_hd__nor2_1 _17011_ (.A(_08152_),
    .B(_08205_),
    .Y(_08206_));
 sky130_fd_sc_hd__nor2_1 _17012_ (.A(_08093_),
    .B(_08148_),
    .Y(_08207_));
 sky130_fd_sc_hd__inv_2 _17013_ (.A(_08207_),
    .Y(_08208_));
 sky130_fd_sc_hd__and3_1 _17014_ (.A(_08152_),
    .B(_08205_),
    .C(_08208_),
    .X(_08209_));
 sky130_fd_sc_hd__a21oi_1 _17015_ (.A1(_08152_),
    .A2(_08208_),
    .B1(_08205_),
    .Y(_08210_));
 sky130_fd_sc_hd__or3_1 _17016_ (.A(net278),
    .B(_08209_),
    .C(_08210_),
    .X(_08211_));
 sky130_fd_sc_hd__a21bo_1 _17017_ (.A1(net354),
    .A2(net273),
    .B1_N(net656),
    .X(_08212_));
 sky130_fd_sc_hd__inv_2 _17018_ (.A(_08212_),
    .Y(_08213_));
 sky130_fd_sc_hd__or3b_1 _17019_ (.A(net656),
    .B(net271),
    .C_N(net354),
    .X(_08214_));
 sky130_fd_sc_hd__o21bai_2 _17020_ (.A1(_08156_),
    .A2(_08159_),
    .B1_N(_08155_),
    .Y(_08216_));
 sky130_fd_sc_hd__a21oi_1 _17021_ (.A1(_08212_),
    .A2(_08214_),
    .B1(_08216_),
    .Y(_08217_));
 sky130_fd_sc_hd__a31o_1 _17022_ (.A1(_08212_),
    .A2(_08214_),
    .A3(_08216_),
    .B1(net229),
    .X(_08218_));
 sky130_fd_sc_hd__nand2_1 _17023_ (.A(_05334_),
    .B(_05764_),
    .Y(_08219_));
 sky130_fd_sc_hd__xor2_1 _17024_ (.A(_05828_),
    .B(_08219_),
    .X(_08220_));
 sky130_fd_sc_hd__a21boi_1 _17025_ (.A1(_01378_),
    .A2(_02564_),
    .B1_N(_01375_),
    .Y(_08221_));
 sky130_fd_sc_hd__o21ai_1 _17026_ (.A1(_02566_),
    .A2(_08221_),
    .B1(net260),
    .Y(_08222_));
 sky130_fd_sc_hd__a21o_2 _17027_ (.A1(_02566_),
    .A2(_08221_),
    .B1(_08222_),
    .X(_08223_));
 sky130_fd_sc_hd__nor2_1 _17028_ (.A(net658),
    .B(_05873_),
    .Y(_08224_));
 sky130_fd_sc_hd__or3_1 _17029_ (.A(net250),
    .B(_05874_),
    .C(_08224_),
    .X(_08225_));
 sky130_fd_sc_hd__a221o_1 _17030_ (.A1(_05764_),
    .A2(net238),
    .B1(net232),
    .B2(net658),
    .C1(net245),
    .X(_08227_));
 sky130_fd_sc_hd__o21ba_1 _17031_ (.A1(_05334_),
    .A2(net235),
    .B1_N(_08227_),
    .X(_08228_));
 sky130_fd_sc_hd__o22a_1 _17032_ (.A1(net211),
    .A2(_05625_),
    .B1(net203),
    .B2(_06796_),
    .X(_08229_));
 sky130_fd_sc_hd__and4_1 _17033_ (.A(_08223_),
    .B(_08225_),
    .C(_08228_),
    .D(_08229_),
    .X(_08230_));
 sky130_fd_sc_hd__o22a_1 _17034_ (.A1(_08217_),
    .A2(_08218_),
    .B1(_08220_),
    .B2(net252),
    .X(_08231_));
 sky130_fd_sc_hd__and3_1 _17035_ (.A(_08211_),
    .B(_08230_),
    .C(_08231_),
    .X(_08232_));
 sky130_fd_sc_hd__a21oi_1 _17036_ (.A1(net656),
    .A2(net246),
    .B1(_08232_),
    .Y(_08703_));
 sky130_fd_sc_hd__nor2_1 _17037_ (.A(_08147_),
    .B(_08201_),
    .Y(_08233_));
 sky130_fd_sc_hd__nor3_2 _17038_ (.A(_06561_),
    .B(_00221_),
    .C(net266),
    .Y(_08234_));
 sky130_fd_sc_hd__o21a_1 _17039_ (.A1(net266),
    .A2(_08234_),
    .B1(_08174_),
    .X(_08235_));
 sky130_fd_sc_hd__nor2_2 _17040_ (.A(_08174_),
    .B(_08234_),
    .Y(_08237_));
 sky130_fd_sc_hd__a211oi_2 _17041_ (.A1(_08613_),
    .A2(_08626_),
    .B1(_08235_),
    .C1(_08237_),
    .Y(_08238_));
 sky130_fd_sc_hd__a21oi_1 _17042_ (.A1(net762),
    .A2(net170),
    .B1(_08238_),
    .Y(_08239_));
 sky130_fd_sc_hd__and3_1 _17043_ (.A(net762),
    .B(net170),
    .C(_08238_),
    .X(_08240_));
 sky130_fd_sc_hd__nor2_1 _17044_ (.A(_08239_),
    .B(_08240_),
    .Y(_08241_));
 sky130_fd_sc_hd__o21a_1 _17045_ (.A1(_08177_),
    .A2(_08184_),
    .B1(_08241_),
    .X(_08242_));
 sky130_fd_sc_hd__nor3_1 _17046_ (.A(_08177_),
    .B(_08184_),
    .C(_08241_),
    .Y(_08243_));
 sky130_fd_sc_hd__nor2_1 _17047_ (.A(_08242_),
    .B(_08243_),
    .Y(_08244_));
 sky130_fd_sc_hd__and2_1 _17048_ (.A(_08180_),
    .B(_08244_),
    .X(_08245_));
 sky130_fd_sc_hd__nor2_1 _17049_ (.A(_08180_),
    .B(_08244_),
    .Y(_08246_));
 sky130_fd_sc_hd__or2_1 _17050_ (.A(_08245_),
    .B(_08246_),
    .X(_08248_));
 sky130_fd_sc_hd__o21ba_1 _17051_ (.A1(_08189_),
    .A2(_08192_),
    .B1_N(_08248_),
    .X(_08249_));
 sky130_fd_sc_hd__or3b_1 _17052_ (.A(_08189_),
    .B(_08192_),
    .C_N(_08248_),
    .X(_08250_));
 sky130_fd_sc_hd__nand2b_2 _17053_ (.A_N(_08249_),
    .B(_08250_),
    .Y(_08251_));
 sky130_fd_sc_hd__nand2_1 _17054_ (.A(_08196_),
    .B(_08200_),
    .Y(_08252_));
 sky130_fd_sc_hd__xor2_1 _17055_ (.A(_08251_),
    .B(_08252_),
    .X(_08253_));
 sky130_fd_sc_hd__and2b_1 _17056_ (.A_N(_08253_),
    .B(_08233_),
    .X(_08254_));
 sky130_fd_sc_hd__and2b_1 _17057_ (.A_N(_08233_),
    .B(_08253_),
    .X(_08255_));
 sky130_fd_sc_hd__nor2_1 _17058_ (.A(_08254_),
    .B(_08255_),
    .Y(_08256_));
 sky130_fd_sc_hd__o22ai_4 _17059_ (.A1(_08201_),
    .A2(_08202_),
    .B1(_08205_),
    .B2(_08208_),
    .Y(_08257_));
 sky130_fd_sc_hd__nor2_1 _17060_ (.A(_08206_),
    .B(_08257_),
    .Y(_08259_));
 sky130_fd_sc_hd__o21a_1 _17061_ (.A1(_08206_),
    .A2(_08257_),
    .B1(_08256_),
    .X(_08260_));
 sky130_fd_sc_hd__xor2_1 _17062_ (.A(_08256_),
    .B(_08259_),
    .X(_08261_));
 sky130_fd_sc_hd__nor2_1 _17063_ (.A(net278),
    .B(_08261_),
    .Y(_08262_));
 sky130_fd_sc_hd__a21bo_2 _17064_ (.A1(net343),
    .A2(net273),
    .B1_N(net646),
    .X(_08263_));
 sky130_fd_sc_hd__or3b_4 _17065_ (.A(net646),
    .B(net271),
    .C_N(net348),
    .X(_08264_));
 sky130_fd_sc_hd__and2_2 _17066_ (.A(_08214_),
    .B(_08216_),
    .X(_08265_));
 sky130_fd_sc_hd__o211ai_4 _17067_ (.A1(_08213_),
    .A2(_08265_),
    .B1(_08264_),
    .C1(_08263_),
    .Y(_08266_));
 sky130_fd_sc_hd__a211o_1 _17068_ (.A1(_08263_),
    .A2(_08264_),
    .B1(_08265_),
    .C1(_08213_),
    .X(_08267_));
 sky130_fd_sc_hd__o211ai_1 _17069_ (.A1(_05408_),
    .A2(_05762_),
    .B1(_05829_),
    .C1(_05334_),
    .Y(_08268_));
 sky130_fd_sc_hd__nor2_1 _17070_ (.A(_02568_),
    .B(net255),
    .Y(_08270_));
 sky130_fd_sc_hd__o21a_2 _17071_ (.A1(_01145_),
    .A2(_02567_),
    .B1(_08270_),
    .X(_08271_));
 sky130_fd_sc_hd__a21oi_1 _17072_ (.A1(net647),
    .A2(_05874_),
    .B1(net250),
    .Y(_08272_));
 sky130_fd_sc_hd__o21a_1 _17073_ (.A1(net647),
    .A2(_05874_),
    .B1(_08272_),
    .X(_08273_));
 sky130_fd_sc_hd__a221o_1 _17074_ (.A1(_05763_),
    .A2(net238),
    .B1(net232),
    .B2(net647),
    .C1(net245),
    .X(_08274_));
 sky130_fd_sc_hd__a21o_1 _17075_ (.A1(_05408_),
    .A2(net236),
    .B1(_08274_),
    .X(_08275_));
 sky130_fd_sc_hd__o32a_1 _17076_ (.A1(net577),
    .A2(_05939_),
    .A3(_06215_),
    .B1(net211),
    .B2(_05658_),
    .X(_08276_));
 sky130_fd_sc_hd__or4b_1 _17077_ (.A(_08271_),
    .B(_08273_),
    .C(_08275_),
    .D_N(_08276_),
    .X(_08277_));
 sky130_fd_sc_hd__a31o_1 _17078_ (.A1(_05830_),
    .A2(_05840_),
    .A3(_08268_),
    .B1(_08277_),
    .X(_08278_));
 sky130_fd_sc_hd__a31o_1 _17079_ (.A1(net230),
    .A2(_08266_),
    .A3(_08267_),
    .B1(_08278_),
    .X(_08279_));
 sky130_fd_sc_hd__o2bb2a_1 _17080_ (.A1_N(net647),
    .A2_N(net246),
    .B1(_08262_),
    .B2(_08279_),
    .X(_08704_));
 sky130_fd_sc_hd__or3b_1 _17081_ (.A(_06561_),
    .B(_06692_),
    .C_N(_00221_),
    .X(_08281_));
 sky130_fd_sc_hd__a32o_1 _17082_ (.A1(net448),
    .A2(net771),
    .A3(_00221_),
    .B1(net458),
    .B2(net758),
    .X(_08282_));
 sky130_fd_sc_hd__and3_2 _17083_ (.A(_06179_),
    .B(_08281_),
    .C(_08282_),
    .X(_08283_));
 sky130_fd_sc_hd__o21ai_2 _17084_ (.A1(_08237_),
    .A2(_08240_),
    .B1(_08283_),
    .Y(_08284_));
 sky130_fd_sc_hd__or3_1 _17085_ (.A(_08237_),
    .B(_08240_),
    .C(_08283_),
    .X(_08285_));
 sky130_fd_sc_hd__and2_1 _17086_ (.A(_08284_),
    .B(_08285_),
    .X(_08286_));
 sky130_fd_sc_hd__o21a_1 _17087_ (.A1(_08242_),
    .A2(_08245_),
    .B1(_08286_),
    .X(_08287_));
 sky130_fd_sc_hd__nor3_1 _17088_ (.A(_08242_),
    .B(_08245_),
    .C(_08286_),
    .Y(_08288_));
 sky130_fd_sc_hd__nor2_2 _17089_ (.A(_08287_),
    .B(_08288_),
    .Y(_08289_));
 sky130_fd_sc_hd__nor2_1 _17090_ (.A(_08196_),
    .B(_08251_),
    .Y(_08291_));
 sky130_fd_sc_hd__or2_1 _17091_ (.A(_08249_),
    .B(_08291_),
    .X(_08292_));
 sky130_fd_sc_hd__xnor2_1 _17092_ (.A(_08289_),
    .B(_08292_),
    .Y(_08293_));
 sky130_fd_sc_hd__nor3_1 _17093_ (.A(_08200_),
    .B(_08251_),
    .C(_08293_),
    .Y(_08294_));
 sky130_fd_sc_hd__o21ai_1 _17094_ (.A1(_08200_),
    .A2(_08251_),
    .B1(_08293_),
    .Y(_08295_));
 sky130_fd_sc_hd__and2b_1 _17095_ (.A_N(_08294_),
    .B(_08295_),
    .X(_08296_));
 sky130_fd_sc_hd__nor3_1 _17096_ (.A(_08254_),
    .B(_08260_),
    .C(_08296_),
    .Y(_08297_));
 sky130_fd_sc_hd__o21a_1 _17097_ (.A1(_08254_),
    .A2(_08260_),
    .B1(_08296_),
    .X(_08298_));
 sky130_fd_sc_hd__a21boi_4 _17098_ (.A1(net336),
    .A2(net273),
    .B1_N(net638),
    .Y(_08299_));
 sky130_fd_sc_hd__inv_2 _17099_ (.A(_08299_),
    .Y(_08300_));
 sky130_fd_sc_hd__and3b_1 _17100_ (.A_N(net638),
    .B(net273),
    .C(net336),
    .X(_08302_));
 sky130_fd_sc_hd__o211a_1 _17101_ (.A1(_08299_),
    .A2(_08302_),
    .B1(_08263_),
    .C1(_08266_),
    .X(_08303_));
 sky130_fd_sc_hd__a211o_1 _17102_ (.A1(_08263_),
    .A2(_08266_),
    .B1(_08299_),
    .C1(_08302_),
    .X(_08304_));
 sky130_fd_sc_hd__or3b_1 _17103_ (.A(net229),
    .B(_08303_),
    .C_N(_08304_),
    .X(_08305_));
 sky130_fd_sc_hd__o211a_1 _17104_ (.A1(_05582_),
    .A2(_05831_),
    .B1(_05830_),
    .C1(_05407_),
    .X(_08306_));
 sky130_fd_sc_hd__nor2_1 _17105_ (.A(_01141_),
    .B(_02568_),
    .Y(_08307_));
 sky130_fd_sc_hd__o21ai_1 _17106_ (.A1(_02570_),
    .A2(_08307_),
    .B1(net260),
    .Y(_08308_));
 sky130_fd_sc_hd__a21o_2 _17107_ (.A1(_02570_),
    .A2(_08307_),
    .B1(_08308_),
    .X(_08309_));
 sky130_fd_sc_hd__a21oi_1 _17108_ (.A1(net646),
    .A2(_05874_),
    .B1(net637),
    .Y(_08310_));
 sky130_fd_sc_hd__or3_1 _17109_ (.A(net250),
    .B(_05875_),
    .C(_08310_),
    .X(_08311_));
 sky130_fd_sc_hd__o2bb2a_1 _17110_ (.A1_N(net637),
    .A2_N(net232),
    .B1(_05942_),
    .B2(_05831_),
    .X(_08313_));
 sky130_fd_sc_hd__o211a_1 _17111_ (.A1(_05583_),
    .A2(_05945_),
    .B1(_08313_),
    .C1(_05880_),
    .X(_08314_));
 sky130_fd_sc_hd__o32a_1 _17112_ (.A1(net569),
    .A2(net203),
    .A3(_06293_),
    .B1(net209),
    .B2(_05699_),
    .X(_08315_));
 sky130_fd_sc_hd__and3_1 _17113_ (.A(_08311_),
    .B(_08314_),
    .C(_08315_),
    .X(_08316_));
 sky130_fd_sc_hd__o311a_1 _17114_ (.A1(_05832_),
    .A2(net252),
    .A3(_08306_),
    .B1(_08309_),
    .C1(_08316_),
    .X(_08317_));
 sky130_fd_sc_hd__o31a_1 _17115_ (.A1(net278),
    .A2(_08297_),
    .A3(_08298_),
    .B1(_08317_),
    .X(_08318_));
 sky130_fd_sc_hd__a22oi_1 _17116_ (.A1(net638),
    .A2(net245),
    .B1(_08305_),
    .B2(_08318_),
    .Y(_08705_));
 sky130_fd_sc_hd__o31a_1 _17117_ (.A1(_08254_),
    .A2(_08260_),
    .A3(_08294_),
    .B1(_08295_),
    .X(_08319_));
 sky130_fd_sc_hd__nand2_1 _17118_ (.A(_08289_),
    .B(_08291_),
    .Y(_08320_));
 sky130_fd_sc_hd__and3_1 _17119_ (.A(net762),
    .B(_08626_),
    .C(_07128_),
    .X(_08321_));
 sky130_fd_sc_hd__o41a_1 _17120_ (.A1(net762),
    .A2(_06561_),
    .A3(_00221_),
    .A4(net266),
    .B1(_08284_),
    .X(_08323_));
 sky130_fd_sc_hd__xnor2_1 _17121_ (.A(_08321_),
    .B(_08323_),
    .Y(_08324_));
 sky130_fd_sc_hd__a21o_1 _17122_ (.A1(_08249_),
    .A2(_08289_),
    .B1(_08287_),
    .X(_08325_));
 sky130_fd_sc_hd__nand2_1 _17123_ (.A(_08324_),
    .B(_08325_),
    .Y(_08326_));
 sky130_fd_sc_hd__or2_1 _17124_ (.A(_08324_),
    .B(_08325_),
    .X(_08327_));
 sky130_fd_sc_hd__nand2_1 _17125_ (.A(_08326_),
    .B(_08327_),
    .Y(_08328_));
 sky130_fd_sc_hd__or2_1 _17126_ (.A(_08320_),
    .B(_08328_),
    .X(_08329_));
 sky130_fd_sc_hd__nand2_1 _17127_ (.A(_08320_),
    .B(_08328_),
    .Y(_08330_));
 sky130_fd_sc_hd__and2_1 _17128_ (.A(_08329_),
    .B(_08330_),
    .X(_08331_));
 sky130_fd_sc_hd__nand2_1 _17129_ (.A(_08319_),
    .B(_08331_),
    .Y(_08332_));
 sky130_fd_sc_hd__or2_1 _17130_ (.A(_08319_),
    .B(_08331_),
    .X(_08334_));
 sky130_fd_sc_hd__and3_1 _17131_ (.A(net280),
    .B(_08332_),
    .C(_08334_),
    .X(_08335_));
 sky130_fd_sc_hd__a21o_1 _17132_ (.A1(net329),
    .A2(net273),
    .B1(_03258_),
    .X(_08336_));
 sky130_fd_sc_hd__inv_2 _17133_ (.A(_08336_),
    .Y(_08337_));
 sky130_fd_sc_hd__and3_1 _17134_ (.A(net329),
    .B(_03258_),
    .C(net273),
    .X(_08338_));
 sky130_fd_sc_hd__o211ai_1 _17135_ (.A1(_08337_),
    .A2(_08338_),
    .B1(_08300_),
    .C1(_08304_),
    .Y(_08339_));
 sky130_fd_sc_hd__a211o_1 _17136_ (.A1(_08300_),
    .A2(_08304_),
    .B1(_08337_),
    .C1(_08338_),
    .X(_08340_));
 sky130_fd_sc_hd__a211o_1 _17137_ (.A1(_05666_),
    .A2(_05833_),
    .B1(_05832_),
    .C1(_05582_),
    .X(_08341_));
 sky130_fd_sc_hd__xnor2_4 _17138_ (.A(_00893_),
    .B(_02571_),
    .Y(_08342_));
 sky130_fd_sc_hd__nor2_1 _17139_ (.A(net628),
    .B(_05875_),
    .Y(_08343_));
 sky130_fd_sc_hd__or3_1 _17140_ (.A(net250),
    .B(_05876_),
    .C(_08343_),
    .X(_08345_));
 sky130_fd_sc_hd__a221o_1 _17141_ (.A1(_05833_),
    .A2(net239),
    .B1(net232),
    .B2(net628),
    .C1(net245),
    .X(_08346_));
 sky130_fd_sc_hd__o21ba_1 _17142_ (.A1(_05666_),
    .A2(_05945_),
    .B1_N(_08346_),
    .X(_08347_));
 sky130_fd_sc_hd__o21a_1 _17143_ (.A1(net208),
    .A2(_05730_),
    .B1(_08347_),
    .X(_08348_));
 sky130_fd_sc_hd__o211a_1 _17144_ (.A1(net203),
    .A2(_07119_),
    .B1(_08345_),
    .C1(_08348_),
    .X(_08349_));
 sky130_fd_sc_hd__o21ai_2 _17145_ (.A1(net257),
    .A2(_08342_),
    .B1(_08349_),
    .Y(_08350_));
 sky130_fd_sc_hd__a31o_1 _17146_ (.A1(_05951_),
    .A2(_08339_),
    .A3(_08340_),
    .B1(_08350_),
    .X(_08351_));
 sky130_fd_sc_hd__a31o_1 _17147_ (.A1(_05835_),
    .A2(_05840_),
    .A3(_08341_),
    .B1(_08351_),
    .X(_08352_));
 sky130_fd_sc_hd__o22a_1 _17148_ (.A1(_03258_),
    .A2(_05880_),
    .B1(_08335_),
    .B2(_08352_),
    .X(_08707_));
 sky130_fd_sc_hd__a211o_1 _17149_ (.A1(_08626_),
    .A2(_08284_),
    .B1(net266),
    .C1(_05001_),
    .X(_08353_));
 sky130_fd_sc_hd__a41o_1 _17150_ (.A1(_08326_),
    .A2(_08329_),
    .A3(_08332_),
    .A4(_08353_),
    .B1(net277),
    .X(_08355_));
 sky130_fd_sc_hd__nand2_1 _17151_ (.A(_05735_),
    .B(_05837_),
    .Y(_08356_));
 sky130_fd_sc_hd__nor2_1 _17152_ (.A(net271),
    .B(_08356_),
    .Y(_08357_));
 sky130_fd_sc_hd__and2_1 _17153_ (.A(net621),
    .B(net271),
    .X(_08358_));
 sky130_fd_sc_hd__a211o_1 _17154_ (.A1(_08336_),
    .A2(_08340_),
    .B1(_08357_),
    .C1(_08358_),
    .X(_08359_));
 sky130_fd_sc_hd__o211a_1 _17155_ (.A1(_08357_),
    .A2(_08358_),
    .B1(_08336_),
    .C1(_08340_),
    .X(_08360_));
 sky130_fd_sc_hd__or3b_1 _17156_ (.A(_08360_),
    .B(_05952_),
    .C_N(_08359_),
    .X(_08361_));
 sky130_fd_sc_hd__a21boi_4 _17157_ (.A1(_00893_),
    .A2(_02571_),
    .B1_N(_00890_),
    .Y(_08362_));
 sky130_fd_sc_hd__a21oi_2 _17158_ (.A1(_02573_),
    .A2(_08362_),
    .B1(net255),
    .Y(_08363_));
 sky130_fd_sc_hd__o21ai_4 _17159_ (.A1(_02573_),
    .A2(_08362_),
    .B1(_08363_),
    .Y(_08364_));
 sky130_fd_sc_hd__a21oi_1 _17160_ (.A1(net620),
    .A2(_05876_),
    .B1(net250),
    .Y(_08366_));
 sky130_fd_sc_hd__o21ai_1 _17161_ (.A1(net620),
    .A2(_05876_),
    .B1(_08366_),
    .Y(_08367_));
 sky130_fd_sc_hd__a221o_1 _17162_ (.A1(_05837_),
    .A2(net238),
    .B1(net232),
    .B2(net620),
    .C1(net245),
    .X(_08368_));
 sky130_fd_sc_hd__o21ba_1 _17163_ (.A1(_05735_),
    .A2(net235),
    .B1_N(_08368_),
    .X(_08369_));
 sky130_fd_sc_hd__or4_1 _17164_ (.A(net568),
    .B(net585),
    .C(net203),
    .D(_06122_),
    .X(_08370_));
 sky130_fd_sc_hd__o211a_1 _17165_ (.A1(net208),
    .A2(_05755_),
    .B1(_08369_),
    .C1(_08370_),
    .X(_08371_));
 sky130_fd_sc_hd__and3_1 _17166_ (.A(_08364_),
    .B(_08367_),
    .C(_08371_),
    .X(_08372_));
 sky130_fd_sc_hd__and3_1 _17167_ (.A(_05666_),
    .B(_05835_),
    .C(_08356_),
    .X(_08373_));
 sky130_fd_sc_hd__a21oi_1 _17168_ (.A1(_05666_),
    .A2(_05835_),
    .B1(_08356_),
    .Y(_08374_));
 sky130_fd_sc_hd__o31a_1 _17169_ (.A1(net252),
    .A2(_08373_),
    .A3(_08374_),
    .B1(_08372_),
    .X(_08375_));
 sky130_fd_sc_hd__a32oi_1 _17170_ (.A1(_08355_),
    .A2(_08361_),
    .A3(_08375_),
    .B1(net245),
    .B2(net621),
    .Y(_08708_));
 sky130_fd_sc_hd__and3b_1 _17171_ (.A_N(net68),
    .B(net67),
    .C(net34),
    .X(_08377_));
 sky130_fd_sc_hd__nand3b_1 _17172_ (.A_N(net68),
    .B(net67),
    .C(net34),
    .Y(_08378_));
 sky130_fd_sc_hd__or3b_2 _17173_ (.A(net26),
    .B(net25),
    .C_N(net23),
    .X(_08379_));
 sky130_fd_sc_hd__or4b_1 _17174_ (.A(net18),
    .B(net21),
    .C(net20),
    .D_N(net22),
    .X(_08380_));
 sky130_fd_sc_hd__or4_1 _17175_ (.A(net14),
    .B(net17),
    .C(net16),
    .D(net19),
    .X(_08381_));
 sky130_fd_sc_hd__or4_1 _17176_ (.A(net32),
    .B(net4),
    .C(net3),
    .D(net6),
    .X(_08382_));
 sky130_fd_sc_hd__or4_1 _17177_ (.A(net29),
    .B(net31),
    .C(net30),
    .D(net33),
    .X(_08383_));
 sky130_fd_sc_hd__or4_1 _17178_ (.A(net5),
    .B(net8),
    .C(net7),
    .D(net10),
    .X(_08384_));
 sky130_fd_sc_hd__or4_1 _17179_ (.A(net9),
    .B(net12),
    .C(net11),
    .D(net15),
    .X(_08385_));
 sky130_fd_sc_hd__or4_2 _17180_ (.A(_08382_),
    .B(_08383_),
    .C(_08384_),
    .D(_08385_),
    .X(_08387_));
 sky130_fd_sc_hd__nor4_2 _17181_ (.A(_08379_),
    .B(_08380_),
    .C(_08381_),
    .D(_08387_),
    .Y(_08388_));
 sky130_fd_sc_hd__and2b_1 _17182_ (.A_N(net28),
    .B(net222),
    .X(_08389_));
 sky130_fd_sc_hd__nor2_8 _17183_ (.A(net13),
    .B(net2),
    .Y(_08390_));
 sky130_fd_sc_hd__nand2_2 _17184_ (.A(net24),
    .B(_08390_),
    .Y(_08391_));
 sky130_fd_sc_hd__and4_2 _17185_ (.A(net24),
    .B(_03313_),
    .C(net1),
    .D(_08390_),
    .X(_08392_));
 sky130_fd_sc_hd__nand2_1 _17186_ (.A(net28),
    .B(net222),
    .Y(_08393_));
 sky130_fd_sc_hd__nor3_1 _17187_ (.A(net27),
    .B(_08391_),
    .C(_08393_),
    .Y(_08394_));
 sky130_fd_sc_hd__or4_1 _17188_ (.A(net14),
    .B(net19),
    .C(net21),
    .D(net20),
    .X(_08395_));
 sky130_fd_sc_hd__or4_1 _17189_ (.A(net29),
    .B(net33),
    .C(net4),
    .D(net3),
    .X(_08396_));
 sky130_fd_sc_hd__or4_1 _17190_ (.A(net8),
    .B(net7),
    .C(net9),
    .D(net15),
    .X(_08398_));
 sky130_fd_sc_hd__or4_1 _17191_ (.A(_08379_),
    .B(_08395_),
    .C(_08396_),
    .D(_08398_),
    .X(_08399_));
 sky130_fd_sc_hd__or4b_1 _17192_ (.A(net17),
    .B(net16),
    .C(net18),
    .D_N(net22),
    .X(_08400_));
 sky130_fd_sc_hd__or4_1 _17193_ (.A(net31),
    .B(net30),
    .C(net32),
    .D(net6),
    .X(_08401_));
 sky130_fd_sc_hd__or4_1 _17194_ (.A(net5),
    .B(net10),
    .C(net12),
    .D(net11),
    .X(_08402_));
 sky130_fd_sc_hd__or3_1 _17195_ (.A(_08400_),
    .B(_08401_),
    .C(_08402_),
    .X(_08403_));
 sky130_fd_sc_hd__or3_4 _17196_ (.A(net28),
    .B(_08399_),
    .C(_08403_),
    .X(_08404_));
 sky130_fd_sc_hd__a221o_1 _17197_ (.A1(_08389_),
    .A2(_08392_),
    .B1(net130),
    .B2(\salida[32] ),
    .C1(net922),
    .X(_08405_));
 sky130_fd_sc_hd__and4b_1 _17198_ (.A_N(net24),
    .B(net27),
    .C(_08389_),
    .D(_08390_),
    .X(_08406_));
 sky130_fd_sc_hd__and2_1 _17199_ (.A(\salida[0] ),
    .B(net123),
    .X(_08407_));
 sky130_fd_sc_hd__o221a_1 _17200_ (.A1(net83),
    .A2(net923),
    .B1(_08405_),
    .B2(_08407_),
    .C1(net934),
    .X(_00004_));
 sky130_fd_sc_hd__a21o_1 _17201_ (.A1(\salida[33] ),
    .A2(net127),
    .B1(net919),
    .X(_08409_));
 sky130_fd_sc_hd__and2_1 _17202_ (.A(\salida[1] ),
    .B(net123),
    .X(_08410_));
 sky130_fd_sc_hd__o221a_1 _17203_ (.A1(net94),
    .A2(net923),
    .B1(_08409_),
    .B2(_08410_),
    .C1(net933),
    .X(_00005_));
 sky130_fd_sc_hd__a21o_1 _17204_ (.A1(\salida[34] ),
    .A2(net127),
    .B1(net919),
    .X(_08411_));
 sky130_fd_sc_hd__and2_1 _17205_ (.A(\salida[2] ),
    .B(net123),
    .X(_08412_));
 sky130_fd_sc_hd__o221a_1 _17206_ (.A1(net105),
    .A2(net923),
    .B1(_08411_),
    .B2(_08412_),
    .C1(net933),
    .X(_00006_));
 sky130_fd_sc_hd__a21o_1 _17207_ (.A1(\salida[35] ),
    .A2(net127),
    .B1(net919),
    .X(_08413_));
 sky130_fd_sc_hd__and2_1 _17208_ (.A(\salida[3] ),
    .B(net123),
    .X(_08414_));
 sky130_fd_sc_hd__o221a_1 _17209_ (.A1(net108),
    .A2(net923),
    .B1(_08413_),
    .B2(_08414_),
    .C1(net933),
    .X(_00007_));
 sky130_fd_sc_hd__a21o_1 _17210_ (.A1(\salida[36] ),
    .A2(net127),
    .B1(net919),
    .X(_08416_));
 sky130_fd_sc_hd__and2_1 _17211_ (.A(\salida[4] ),
    .B(net123),
    .X(_08417_));
 sky130_fd_sc_hd__o221a_1 _17212_ (.A1(net109),
    .A2(net923),
    .B1(_08416_),
    .B2(_08417_),
    .C1(net934),
    .X(_00008_));
 sky130_fd_sc_hd__a21o_1 _17213_ (.A1(\salida[37] ),
    .A2(net130),
    .B1(net922),
    .X(_08418_));
 sky130_fd_sc_hd__and2_1 _17214_ (.A(\salida[5] ),
    .B(net126),
    .X(_08419_));
 sky130_fd_sc_hd__o221a_1 _17215_ (.A1(net110),
    .A2(net926),
    .B1(_08418_),
    .B2(_08419_),
    .C1(net934),
    .X(_00009_));
 sky130_fd_sc_hd__a21o_1 _17216_ (.A1(\salida[38] ),
    .A2(net127),
    .B1(net919),
    .X(_08420_));
 sky130_fd_sc_hd__and2_1 _17217_ (.A(\salida[6] ),
    .B(net123),
    .X(_08421_));
 sky130_fd_sc_hd__o221a_1 _17218_ (.A1(net111),
    .A2(net923),
    .B1(_08420_),
    .B2(_08421_),
    .C1(net934),
    .X(_00010_));
 sky130_fd_sc_hd__a21o_1 _17219_ (.A1(\salida[39] ),
    .A2(net127),
    .B1(net919),
    .X(_08422_));
 sky130_fd_sc_hd__and2_1 _17220_ (.A(\salida[7] ),
    .B(net123),
    .X(_08424_));
 sky130_fd_sc_hd__o221a_1 _17221_ (.A1(net112),
    .A2(net923),
    .B1(_08422_),
    .B2(_08424_),
    .C1(net935),
    .X(_00011_));
 sky130_fd_sc_hd__a21o_1 _17222_ (.A1(\salida[40] ),
    .A2(net127),
    .B1(net919),
    .X(_08425_));
 sky130_fd_sc_hd__and2_1 _17223_ (.A(\salida[8] ),
    .B(net123),
    .X(_08426_));
 sky130_fd_sc_hd__o221a_1 _17224_ (.A1(net113),
    .A2(net923),
    .B1(_08425_),
    .B2(_08426_),
    .C1(net934),
    .X(_00012_));
 sky130_fd_sc_hd__a21o_1 _17225_ (.A1(\salida[41] ),
    .A2(net127),
    .B1(net919),
    .X(_08427_));
 sky130_fd_sc_hd__and2_1 _17226_ (.A(\salida[9] ),
    .B(net123),
    .X(_08428_));
 sky130_fd_sc_hd__o221a_1 _17227_ (.A1(net114),
    .A2(net923),
    .B1(_08427_),
    .B2(_08428_),
    .C1(net933),
    .X(_00013_));
 sky130_fd_sc_hd__a21o_1 _17228_ (.A1(\salida[42] ),
    .A2(net127),
    .B1(net919),
    .X(_08429_));
 sky130_fd_sc_hd__and2_1 _17229_ (.A(\salida[10] ),
    .B(net126),
    .X(_08430_));
 sky130_fd_sc_hd__o221a_1 _17230_ (.A1(net84),
    .A2(net926),
    .B1(_08429_),
    .B2(_08430_),
    .C1(net935),
    .X(_00014_));
 sky130_fd_sc_hd__a21o_1 _17231_ (.A1(\salida[43] ),
    .A2(net129),
    .B1(net921),
    .X(_08432_));
 sky130_fd_sc_hd__and2_1 _17232_ (.A(\salida[11] ),
    .B(net125),
    .X(_08433_));
 sky130_fd_sc_hd__o221a_1 _17233_ (.A1(net85),
    .A2(net925),
    .B1(_08432_),
    .B2(_08433_),
    .C1(net937),
    .X(_00015_));
 sky130_fd_sc_hd__a21o_1 _17234_ (.A1(\salida[44] ),
    .A2(net129),
    .B1(net921),
    .X(_08434_));
 sky130_fd_sc_hd__and2_1 _17235_ (.A(\salida[12] ),
    .B(net125),
    .X(_08435_));
 sky130_fd_sc_hd__o221a_1 _17236_ (.A1(net86),
    .A2(net925),
    .B1(_08434_),
    .B2(_08435_),
    .C1(net937),
    .X(_00016_));
 sky130_fd_sc_hd__a21o_1 _17237_ (.A1(\salida[45] ),
    .A2(net127),
    .B1(net919),
    .X(_08436_));
 sky130_fd_sc_hd__and2_1 _17238_ (.A(\salida[13] ),
    .B(net123),
    .X(_08437_));
 sky130_fd_sc_hd__o221a_1 _17239_ (.A1(net87),
    .A2(net923),
    .B1(_08436_),
    .B2(_08437_),
    .C1(net934),
    .X(_00017_));
 sky130_fd_sc_hd__a21o_1 _17240_ (.A1(\salida[46] ),
    .A2(net129),
    .B1(net921),
    .X(_08439_));
 sky130_fd_sc_hd__and2_1 _17241_ (.A(\salida[14] ),
    .B(net125),
    .X(_08440_));
 sky130_fd_sc_hd__o221a_1 _17242_ (.A1(net88),
    .A2(net925),
    .B1(_08439_),
    .B2(_08440_),
    .C1(net937),
    .X(_00018_));
 sky130_fd_sc_hd__a21o_1 _17243_ (.A1(\salida[47] ),
    .A2(net129),
    .B1(net921),
    .X(_08441_));
 sky130_fd_sc_hd__and2_1 _17244_ (.A(\salida[15] ),
    .B(net125),
    .X(_08442_));
 sky130_fd_sc_hd__o221a_1 _17245_ (.A1(net89),
    .A2(net925),
    .B1(_08441_),
    .B2(_08442_),
    .C1(net937),
    .X(_00019_));
 sky130_fd_sc_hd__a21o_1 _17246_ (.A1(\salida[48] ),
    .A2(net128),
    .B1(net920),
    .X(_08443_));
 sky130_fd_sc_hd__and2_1 _17247_ (.A(\salida[16] ),
    .B(net125),
    .X(_08444_));
 sky130_fd_sc_hd__o221a_1 _17248_ (.A1(net90),
    .A2(net924),
    .B1(_08443_),
    .B2(_08444_),
    .C1(net936),
    .X(_00020_));
 sky130_fd_sc_hd__a21o_1 _17249_ (.A1(\salida[49] ),
    .A2(net128),
    .B1(net920),
    .X(_08445_));
 sky130_fd_sc_hd__and2_1 _17250_ (.A(\salida[17] ),
    .B(net124),
    .X(_08447_));
 sky130_fd_sc_hd__o221a_1 _17251_ (.A1(net91),
    .A2(net924),
    .B1(_08445_),
    .B2(_08447_),
    .C1(net936),
    .X(_00021_));
 sky130_fd_sc_hd__a21o_1 _17252_ (.A1(\salida[50] ),
    .A2(net128),
    .B1(net920),
    .X(_08448_));
 sky130_fd_sc_hd__and2_1 _17253_ (.A(\salida[18] ),
    .B(net124),
    .X(_08449_));
 sky130_fd_sc_hd__o221a_1 _17254_ (.A1(net92),
    .A2(net924),
    .B1(_08448_),
    .B2(_08449_),
    .C1(net937),
    .X(_00022_));
 sky130_fd_sc_hd__a21o_1 _17255_ (.A1(\salida[51] ),
    .A2(net128),
    .B1(net920),
    .X(_08450_));
 sky130_fd_sc_hd__and2_1 _17256_ (.A(\salida[19] ),
    .B(net124),
    .X(_08451_));
 sky130_fd_sc_hd__o221a_1 _17257_ (.A1(net93),
    .A2(net924),
    .B1(_08450_),
    .B2(_08451_),
    .C1(net937),
    .X(_00023_));
 sky130_fd_sc_hd__a21o_1 _17258_ (.A1(\salida[52] ),
    .A2(net128),
    .B1(net920),
    .X(_08452_));
 sky130_fd_sc_hd__and2_1 _17259_ (.A(\salida[20] ),
    .B(net126),
    .X(_08453_));
 sky130_fd_sc_hd__o221a_1 _17260_ (.A1(net95),
    .A2(net924),
    .B1(_08452_),
    .B2(_08453_),
    .C1(net936),
    .X(_00024_));
 sky130_fd_sc_hd__a21o_1 _17261_ (.A1(\salida[53] ),
    .A2(net128),
    .B1(net920),
    .X(_08455_));
 sky130_fd_sc_hd__and2_1 _17262_ (.A(\salida[21] ),
    .B(net125),
    .X(_08456_));
 sky130_fd_sc_hd__o221a_1 _17263_ (.A1(net96),
    .A2(net926),
    .B1(_08455_),
    .B2(_08456_),
    .C1(net936),
    .X(_00025_));
 sky130_fd_sc_hd__a21o_1 _17264_ (.A1(\salida[54] ),
    .A2(net130),
    .B1(net922),
    .X(_08457_));
 sky130_fd_sc_hd__and2_1 _17265_ (.A(\salida[22] ),
    .B(net125),
    .X(_08458_));
 sky130_fd_sc_hd__o221a_1 _17266_ (.A1(net97),
    .A2(net925),
    .B1(_08457_),
    .B2(_08458_),
    .C1(net936),
    .X(_00026_));
 sky130_fd_sc_hd__a21o_1 _17267_ (.A1(\salida[55] ),
    .A2(net128),
    .B1(net920),
    .X(_08459_));
 sky130_fd_sc_hd__and2_1 _17268_ (.A(\salida[23] ),
    .B(net124),
    .X(_08460_));
 sky130_fd_sc_hd__o221a_1 _17269_ (.A1(net98),
    .A2(net924),
    .B1(_08459_),
    .B2(_08460_),
    .C1(net936),
    .X(_00027_));
 sky130_fd_sc_hd__a21o_1 _17270_ (.A1(\salida[56] ),
    .A2(net128),
    .B1(net920),
    .X(_08462_));
 sky130_fd_sc_hd__and2_1 _17271_ (.A(\salida[24] ),
    .B(net124),
    .X(_08463_));
 sky130_fd_sc_hd__o221a_1 _17272_ (.A1(net99),
    .A2(net925),
    .B1(_08462_),
    .B2(_08463_),
    .C1(net936),
    .X(_00028_));
 sky130_fd_sc_hd__a21o_1 _17273_ (.A1(\salida[57] ),
    .A2(net129),
    .B1(net921),
    .X(_08464_));
 sky130_fd_sc_hd__and2_1 _17274_ (.A(\salida[25] ),
    .B(net124),
    .X(_08465_));
 sky130_fd_sc_hd__o221a_1 _17275_ (.A1(net100),
    .A2(net924),
    .B1(_08464_),
    .B2(_08465_),
    .C1(net936),
    .X(_00029_));
 sky130_fd_sc_hd__a21o_1 _17276_ (.A1(\salida[58] ),
    .A2(net128),
    .B1(net920),
    .X(_08466_));
 sky130_fd_sc_hd__and2_1 _17277_ (.A(\salida[26] ),
    .B(net124),
    .X(_08467_));
 sky130_fd_sc_hd__o221a_1 _17278_ (.A1(net101),
    .A2(net924),
    .B1(_08466_),
    .B2(_08467_),
    .C1(net937),
    .X(_00030_));
 sky130_fd_sc_hd__a21o_1 _17279_ (.A1(\salida[59] ),
    .A2(net128),
    .B1(net920),
    .X(_08468_));
 sky130_fd_sc_hd__and2_1 _17280_ (.A(\salida[27] ),
    .B(net124),
    .X(_08470_));
 sky130_fd_sc_hd__o221a_1 _17281_ (.A1(net102),
    .A2(net924),
    .B1(_08468_),
    .B2(_08470_),
    .C1(net938),
    .X(_00031_));
 sky130_fd_sc_hd__a21o_1 _17282_ (.A1(\salida[60] ),
    .A2(net129),
    .B1(net921),
    .X(_08471_));
 sky130_fd_sc_hd__and2_1 _17283_ (.A(\salida[28] ),
    .B(net124),
    .X(_08472_));
 sky130_fd_sc_hd__o221a_1 _17284_ (.A1(net103),
    .A2(net925),
    .B1(_08471_),
    .B2(_08472_),
    .C1(net936),
    .X(_00032_));
 sky130_fd_sc_hd__a21o_1 _17285_ (.A1(\salida[61] ),
    .A2(net129),
    .B1(net921),
    .X(_08473_));
 sky130_fd_sc_hd__and2_1 _17286_ (.A(\salida[29] ),
    .B(net125),
    .X(_08474_));
 sky130_fd_sc_hd__o221a_1 _17287_ (.A1(net104),
    .A2(net925),
    .B1(_08473_),
    .B2(_08474_),
    .C1(net937),
    .X(_00033_));
 sky130_fd_sc_hd__a21o_1 _17288_ (.A1(\salida[62] ),
    .A2(net129),
    .B1(net921),
    .X(_08475_));
 sky130_fd_sc_hd__and2_1 _17289_ (.A(\salida[30] ),
    .B(net125),
    .X(_08476_));
 sky130_fd_sc_hd__o221a_1 _17290_ (.A1(net106),
    .A2(net925),
    .B1(_08475_),
    .B2(_08476_),
    .C1(net937),
    .X(_00034_));
 sky130_fd_sc_hd__a21o_1 _17291_ (.A1(\salida[63] ),
    .A2(net129),
    .B1(net921),
    .X(_08478_));
 sky130_fd_sc_hd__and2_1 _17292_ (.A(\salida[31] ),
    .B(net124),
    .X(_08479_));
 sky130_fd_sc_hd__o221a_2 _17293_ (.A1(net107),
    .A2(net924),
    .B1(_08478_),
    .B2(_08479_),
    .C1(net936),
    .X(_00035_));
 sky130_fd_sc_hd__nand3_4 _17294_ (.A(net34),
    .B(net67),
    .C(net68),
    .Y(_08480_));
 sky130_fd_sc_hd__or4b_4 _17295_ (.A(net24),
    .B(_08480_),
    .C(net27),
    .D_N(_08390_),
    .X(_08481_));
 sky130_fd_sc_hd__nor2_2 _17296_ (.A(net221),
    .B(net265),
    .Y(_08482_));
 sky130_fd_sc_hd__or3_1 _17297_ (.A(net35),
    .B(net219),
    .C(net263),
    .X(_08483_));
 sky130_fd_sc_hd__o211a_1 _17298_ (.A1(net912),
    .A2(net164),
    .B1(_08483_),
    .C1(net929),
    .X(_00036_));
 sky130_fd_sc_hd__or3_1 _17299_ (.A(net46),
    .B(net219),
    .C(net263),
    .X(_08484_));
 sky130_fd_sc_hd__o211a_1 _17300_ (.A1(net902),
    .A2(net165),
    .B1(_08484_),
    .C1(net929),
    .X(_00037_));
 sky130_fd_sc_hd__or3_1 _17301_ (.A(net57),
    .B(net221),
    .C(net265),
    .X(_08486_));
 sky130_fd_sc_hd__o211a_1 _17302_ (.A1(net900),
    .A2(net167),
    .B1(_08486_),
    .C1(net935),
    .X(_00038_));
 sky130_fd_sc_hd__or3_1 _17303_ (.A(net60),
    .B(net221),
    .C(net265),
    .X(_08487_));
 sky130_fd_sc_hd__o211a_1 _17304_ (.A1(net891),
    .A2(net167),
    .B1(_08487_),
    .C1(net935),
    .X(_00039_));
 sky130_fd_sc_hd__or3_1 _17305_ (.A(net61),
    .B(net219),
    .C(net263),
    .X(_08488_));
 sky130_fd_sc_hd__o211a_1 _17306_ (.A1(net879),
    .A2(net165),
    .B1(_08488_),
    .C1(net929),
    .X(_00040_));
 sky130_fd_sc_hd__or3_1 _17307_ (.A(net62),
    .B(net218),
    .C(net262),
    .X(_08489_));
 sky130_fd_sc_hd__o211a_1 _17308_ (.A1(net862),
    .A2(net164),
    .B1(_08489_),
    .C1(net927),
    .X(_00041_));
 sky130_fd_sc_hd__or3_1 _17309_ (.A(net63),
    .B(net219),
    .C(net263),
    .X(_08490_));
 sky130_fd_sc_hd__o211a_1 _17310_ (.A1(\ApproximateM_inst.lob_16.lob1.genblk1[6].genblk1.mux.sel ),
    .A2(net164),
    .B1(_08490_),
    .C1(net929),
    .X(_00042_));
 sky130_fd_sc_hd__or3_1 _17311_ (.A(net64),
    .B(net219),
    .C(net263),
    .X(_08492_));
 sky130_fd_sc_hd__o211a_1 _17312_ (.A1(net841),
    .A2(net165),
    .B1(_08492_),
    .C1(net933),
    .X(_00043_));
 sky130_fd_sc_hd__or3_1 _17313_ (.A(net65),
    .B(net218),
    .C(net262),
    .X(_08493_));
 sky130_fd_sc_hd__o211a_1 _17314_ (.A1(net831),
    .A2(net164),
    .B1(_08493_),
    .C1(net928),
    .X(_00044_));
 sky130_fd_sc_hd__or3_1 _17315_ (.A(net66),
    .B(net220),
    .C(net262),
    .X(_08494_));
 sky130_fd_sc_hd__o211a_1 _17316_ (.A1(net823),
    .A2(net164),
    .B1(_08494_),
    .C1(net928),
    .X(_00045_));
 sky130_fd_sc_hd__or3_1 _17317_ (.A(net36),
    .B(net218),
    .C(net262),
    .X(_08495_));
 sky130_fd_sc_hd__o211a_1 _17318_ (.A1(net812),
    .A2(net164),
    .B1(_08495_),
    .C1(net927),
    .X(_00046_));
 sky130_fd_sc_hd__or3_1 _17319_ (.A(net37),
    .B(net218),
    .C(net262),
    .X(_08496_));
 sky130_fd_sc_hd__o211a_1 _17320_ (.A1(net802),
    .A2(net164),
    .B1(_08496_),
    .C1(net927),
    .X(_00047_));
 sky130_fd_sc_hd__or3_1 _17321_ (.A(net38),
    .B(net218),
    .C(net262),
    .X(_08498_));
 sky130_fd_sc_hd__o211a_1 _17322_ (.A1(net795),
    .A2(net165),
    .B1(_08498_),
    .C1(net929),
    .X(_00048_));
 sky130_fd_sc_hd__or3_1 _17323_ (.A(net39),
    .B(net218),
    .C(net262),
    .X(_08499_));
 sky130_fd_sc_hd__o211a_1 _17324_ (.A1(net779),
    .A2(net164),
    .B1(_08499_),
    .C1(net927),
    .X(_00049_));
 sky130_fd_sc_hd__or3_1 _17325_ (.A(net40),
    .B(net218),
    .C(net262),
    .X(_08500_));
 sky130_fd_sc_hd__o211a_1 _17326_ (.A1(net766),
    .A2(net164),
    .B1(_08500_),
    .C1(net928),
    .X(_00050_));
 sky130_fd_sc_hd__or3_1 _17327_ (.A(net41),
    .B(net219),
    .C(net263),
    .X(_08501_));
 sky130_fd_sc_hd__o211a_1 _17328_ (.A1(net756),
    .A2(net165),
    .B1(_08501_),
    .C1(net929),
    .X(_00051_));
 sky130_fd_sc_hd__or3_1 _17329_ (.A(net42),
    .B(net218),
    .C(net262),
    .X(_08502_));
 sky130_fd_sc_hd__o211a_1 _17330_ (.A1(net747),
    .A2(net164),
    .B1(_08502_),
    .C1(net928),
    .X(_00052_));
 sky130_fd_sc_hd__or3_1 _17331_ (.A(net43),
    .B(net218),
    .C(net263),
    .X(_08504_));
 sky130_fd_sc_hd__o211a_1 _17332_ (.A1(net739),
    .A2(net165),
    .B1(_08504_),
    .C1(net930),
    .X(_00053_));
 sky130_fd_sc_hd__or3_1 _17333_ (.A(net44),
    .B(net218),
    .C(net262),
    .X(_08505_));
 sky130_fd_sc_hd__o211a_1 _17334_ (.A1(net730),
    .A2(net165),
    .B1(_08505_),
    .C1(net929),
    .X(_00054_));
 sky130_fd_sc_hd__or3_1 _17335_ (.A(net45),
    .B(net221),
    .C(net264),
    .X(_08506_));
 sky130_fd_sc_hd__o211a_1 _17336_ (.A1(net721),
    .A2(net167),
    .B1(_08506_),
    .C1(net932),
    .X(_00055_));
 sky130_fd_sc_hd__or3_1 _17337_ (.A(net47),
    .B(net221),
    .C(net265),
    .X(_08507_));
 sky130_fd_sc_hd__o211a_1 _17338_ (.A1(net712),
    .A2(net167),
    .B1(_08507_),
    .C1(net935),
    .X(_00056_));
 sky130_fd_sc_hd__or3_1 _17339_ (.A(net48),
    .B(net220),
    .C(net264),
    .X(_08508_));
 sky130_fd_sc_hd__o211a_1 _17340_ (.A1(net703),
    .A2(net166),
    .B1(_08508_),
    .C1(net931),
    .X(_00057_));
 sky130_fd_sc_hd__or3_1 _17341_ (.A(net49),
    .B(net220),
    .C(net264),
    .X(_08510_));
 sky130_fd_sc_hd__o211a_1 _17342_ (.A1(net695),
    .A2(net166),
    .B1(_08510_),
    .C1(net931),
    .X(_00058_));
 sky130_fd_sc_hd__or3_1 _17343_ (.A(net50),
    .B(net220),
    .C(net264),
    .X(_08511_));
 sky130_fd_sc_hd__o211a_1 _17344_ (.A1(net689),
    .A2(net166),
    .B1(_08511_),
    .C1(net932),
    .X(_00059_));
 sky130_fd_sc_hd__or3_1 _17345_ (.A(net51),
    .B(net220),
    .C(net264),
    .X(_08512_));
 sky130_fd_sc_hd__o211a_1 _17346_ (.A1(net684),
    .A2(net166),
    .B1(_08512_),
    .C1(net931),
    .X(_00060_));
 sky130_fd_sc_hd__or3_1 _17347_ (.A(net52),
    .B(net221),
    .C(net265),
    .X(_08513_));
 sky130_fd_sc_hd__o211a_1 _17348_ (.A1(net671),
    .A2(net167),
    .B1(_08513_),
    .C1(net932),
    .X(_00061_));
 sky130_fd_sc_hd__or3_1 _17349_ (.A(net53),
    .B(net221),
    .C(net265),
    .X(_08514_));
 sky130_fd_sc_hd__o211a_1 _17350_ (.A1(net663),
    .A2(net166),
    .B1(_08514_),
    .C1(net934),
    .X(_00062_));
 sky130_fd_sc_hd__or3_1 _17351_ (.A(net54),
    .B(net220),
    .C(net264),
    .X(_08516_));
 sky130_fd_sc_hd__o211a_1 _17352_ (.A1(net655),
    .A2(net166),
    .B1(_08516_),
    .C1(net932),
    .X(_00063_));
 sky130_fd_sc_hd__or3_1 _17353_ (.A(net55),
    .B(net220),
    .C(net264),
    .X(_08517_));
 sky130_fd_sc_hd__o211a_1 _17354_ (.A1(net645),
    .A2(net166),
    .B1(_08517_),
    .C1(net932),
    .X(_00064_));
 sky130_fd_sc_hd__or3_1 _17355_ (.A(net56),
    .B(net220),
    .C(net264),
    .X(_08518_));
 sky130_fd_sc_hd__o211a_1 _17356_ (.A1(net635),
    .A2(net166),
    .B1(_08518_),
    .C1(net931),
    .X(_00065_));
 sky130_fd_sc_hd__or3_1 _17357_ (.A(net58),
    .B(net220),
    .C(net264),
    .X(_08519_));
 sky130_fd_sc_hd__o211a_1 _17358_ (.A1(net627),
    .A2(net166),
    .B1(_08519_),
    .C1(net931),
    .X(_00066_));
 sky130_fd_sc_hd__or3_1 _17359_ (.A(net59),
    .B(net220),
    .C(net264),
    .X(_08520_));
 sky130_fd_sc_hd__o211a_1 _17360_ (.A1(net619),
    .A2(net166),
    .B1(_08520_),
    .C1(net931),
    .X(_00067_));
 sky130_fd_sc_hd__nor4_4 _17361_ (.A(_03313_),
    .B(_08391_),
    .C(net219),
    .D(_08480_),
    .Y(_08522_));
 sky130_fd_sc_hd__or4_4 _17362_ (.A(_03313_),
    .B(_08391_),
    .C(net219),
    .D(_08480_),
    .X(_08523_));
 sky130_fd_sc_hd__nand2_1 _17363_ (.A(net285),
    .B(net158),
    .Y(_08524_));
 sky130_fd_sc_hd__o211a_1 _17364_ (.A1(net35),
    .A2(net158),
    .B1(_08524_),
    .C1(net933),
    .X(_00068_));
 sky130_fd_sc_hd__nand2_1 _17365_ (.A(net288),
    .B(net158),
    .Y(_08525_));
 sky130_fd_sc_hd__o211a_1 _17366_ (.A1(net46),
    .A2(net158),
    .B1(_08525_),
    .C1(net933),
    .X(_00069_));
 sky130_fd_sc_hd__nand2_1 _17367_ (.A(net295),
    .B(net159),
    .Y(_08526_));
 sky130_fd_sc_hd__o211a_1 _17368_ (.A1(net57),
    .A2(net158),
    .B1(_08526_),
    .C1(net934),
    .X(_00070_));
 sky130_fd_sc_hd__nand2_1 _17369_ (.A(net300),
    .B(net158),
    .Y(_08527_));
 sky130_fd_sc_hd__o211a_1 _17370_ (.A1(net60),
    .A2(net158),
    .B1(_08527_),
    .C1(net934),
    .X(_00071_));
 sky130_fd_sc_hd__nand2_1 _17371_ (.A(net307),
    .B(net158),
    .Y(_08529_));
 sky130_fd_sc_hd__o211a_1 _17372_ (.A1(net61),
    .A2(net158),
    .B1(_08529_),
    .C1(net933),
    .X(_00072_));
 sky130_fd_sc_hd__or2_1 _17373_ (.A(net549),
    .B(net161),
    .X(_08530_));
 sky130_fd_sc_hd__o211a_1 _17374_ (.A1(net62),
    .A2(net156),
    .B1(_08530_),
    .C1(net927),
    .X(_00073_));
 sky130_fd_sc_hd__or2_1 _17375_ (.A(net528),
    .B(net162),
    .X(_08531_));
 sky130_fd_sc_hd__o211a_1 _17376_ (.A1(net63),
    .A2(net156),
    .B1(_08531_),
    .C1(net929),
    .X(_00074_));
 sky130_fd_sc_hd__nand2_1 _17377_ (.A(_03182_),
    .B(net159),
    .Y(_08532_));
 sky130_fd_sc_hd__o211a_1 _17378_ (.A1(net64),
    .A2(net158),
    .B1(_08532_),
    .C1(net933),
    .X(_00075_));
 sky130_fd_sc_hd__or2_1 _17379_ (.A(net511),
    .B(net161),
    .X(_08533_));
 sky130_fd_sc_hd__o211a_1 _17380_ (.A1(net65),
    .A2(net157),
    .B1(_08533_),
    .C1(net928),
    .X(_00076_));
 sky130_fd_sc_hd__or2_1 _17381_ (.A(net503),
    .B(net161),
    .X(_08535_));
 sky130_fd_sc_hd__o211a_1 _17382_ (.A1(net66),
    .A2(net157),
    .B1(_08535_),
    .C1(net928),
    .X(_00077_));
 sky130_fd_sc_hd__or2_1 _17383_ (.A(net494),
    .B(net161),
    .X(_08536_));
 sky130_fd_sc_hd__o211a_1 _17384_ (.A1(net36),
    .A2(net156),
    .B1(_08536_),
    .C1(net927),
    .X(_00078_));
 sky130_fd_sc_hd__or2_1 _17385_ (.A(net484),
    .B(net161),
    .X(_08537_));
 sky130_fd_sc_hd__o211a_1 _17386_ (.A1(net37),
    .A2(net156),
    .B1(_08537_),
    .C1(net927),
    .X(_00079_));
 sky130_fd_sc_hd__or2_1 _17387_ (.A(net479),
    .B(net162),
    .X(_08538_));
 sky130_fd_sc_hd__o211a_1 _17388_ (.A1(net38),
    .A2(net156),
    .B1(_08538_),
    .C1(net927),
    .X(_00080_));
 sky130_fd_sc_hd__or2_1 _17389_ (.A(net472),
    .B(net161),
    .X(_08539_));
 sky130_fd_sc_hd__o211a_1 _17390_ (.A1(net39),
    .A2(net156),
    .B1(_08539_),
    .C1(net927),
    .X(_00081_));
 sky130_fd_sc_hd__or2_1 _17391_ (.A(net462),
    .B(net161),
    .X(_08541_));
 sky130_fd_sc_hd__o211a_1 _17392_ (.A1(net40),
    .A2(net157),
    .B1(_08541_),
    .C1(net928),
    .X(_00082_));
 sky130_fd_sc_hd__or2_1 _17393_ (.A(net450),
    .B(net162),
    .X(_08542_));
 sky130_fd_sc_hd__o211a_1 _17394_ (.A1(net41),
    .A2(net156),
    .B1(_08542_),
    .C1(net929),
    .X(_00083_));
 sky130_fd_sc_hd__or2_1 _17395_ (.A(net444),
    .B(net162),
    .X(_08543_));
 sky130_fd_sc_hd__o211a_1 _17396_ (.A1(net42),
    .A2(net156),
    .B1(_08543_),
    .C1(net927),
    .X(_00084_));
 sky130_fd_sc_hd__or2_1 _17397_ (.A(net433),
    .B(net162),
    .X(_08544_));
 sky130_fd_sc_hd__o211a_1 _17398_ (.A1(net43),
    .A2(net157),
    .B1(_08544_),
    .C1(net930),
    .X(_00085_));
 sky130_fd_sc_hd__or2_1 _17399_ (.A(net426),
    .B(net161),
    .X(_08545_));
 sky130_fd_sc_hd__o211a_1 _17400_ (.A1(net44),
    .A2(net156),
    .B1(_08545_),
    .C1(net930),
    .X(_00086_));
 sky130_fd_sc_hd__or2_1 _17401_ (.A(net417),
    .B(net162),
    .X(_08547_));
 sky130_fd_sc_hd__o211a_1 _17402_ (.A1(net45),
    .A2(net157),
    .B1(_08547_),
    .C1(net929),
    .X(_00087_));
 sky130_fd_sc_hd__or2_1 _17403_ (.A(net410),
    .B(net161),
    .X(_08548_));
 sky130_fd_sc_hd__o211a_1 _17404_ (.A1(net47),
    .A2(net156),
    .B1(_08548_),
    .C1(net930),
    .X(_00088_));
 sky130_fd_sc_hd__or2_1 _17405_ (.A(net401),
    .B(net161),
    .X(_08549_));
 sky130_fd_sc_hd__o211a_1 _17406_ (.A1(net48),
    .A2(net160),
    .B1(_08549_),
    .C1(net931),
    .X(_00089_));
 sky130_fd_sc_hd__or2_1 _17407_ (.A(net393),
    .B(net163),
    .X(_08550_));
 sky130_fd_sc_hd__o211a_1 _17408_ (.A1(net49),
    .A2(net160),
    .B1(_08550_),
    .C1(net931),
    .X(_00090_));
 sky130_fd_sc_hd__or2_1 _17409_ (.A(net384),
    .B(net163),
    .X(_08551_));
 sky130_fd_sc_hd__o211a_1 _17410_ (.A1(net50),
    .A2(net160),
    .B1(_08551_),
    .C1(net932),
    .X(_00091_));
 sky130_fd_sc_hd__or2_1 _17411_ (.A(net376),
    .B(net163),
    .X(_08553_));
 sky130_fd_sc_hd__o211a_1 _17412_ (.A1(net51),
    .A2(net160),
    .B1(_08553_),
    .C1(net931),
    .X(_00092_));
 sky130_fd_sc_hd__or2_1 _17413_ (.A(net367),
    .B(net163),
    .X(_08554_));
 sky130_fd_sc_hd__o211a_1 _17414_ (.A1(net52),
    .A2(net160),
    .B1(_08554_),
    .C1(net932),
    .X(_00093_));
 sky130_fd_sc_hd__or2_1 _17415_ (.A(net359),
    .B(net163),
    .X(_08555_));
 sky130_fd_sc_hd__o211a_1 _17416_ (.A1(net53),
    .A2(_08523_),
    .B1(_08555_),
    .C1(net932),
    .X(_00094_));
 sky130_fd_sc_hd__or2_1 _17417_ (.A(net352),
    .B(net163),
    .X(_08556_));
 sky130_fd_sc_hd__o211a_1 _17418_ (.A1(net54),
    .A2(net160),
    .B1(_08556_),
    .C1(net931),
    .X(_00095_));
 sky130_fd_sc_hd__or2_1 _17419_ (.A(net344),
    .B(net163),
    .X(_08557_));
 sky130_fd_sc_hd__o211a_1 _17420_ (.A1(net55),
    .A2(net160),
    .B1(_08557_),
    .C1(net932),
    .X(_00096_));
 sky130_fd_sc_hd__or2_1 _17421_ (.A(net337),
    .B(net163),
    .X(_08559_));
 sky130_fd_sc_hd__o211a_1 _17422_ (.A1(net56),
    .A2(net160),
    .B1(_08559_),
    .C1(net938),
    .X(_00097_));
 sky130_fd_sc_hd__or2_1 _17423_ (.A(net328),
    .B(_08522_),
    .X(_08560_));
 sky130_fd_sc_hd__o211a_1 _17424_ (.A1(net58),
    .A2(net160),
    .B1(_08560_),
    .C1(net938),
    .X(_00098_));
 sky130_fd_sc_hd__or2_1 _17425_ (.A(net318),
    .B(_08522_),
    .X(_08561_));
 sky130_fd_sc_hd__o211a_1 _17426_ (.A1(net59),
    .A2(net160),
    .B1(_08561_),
    .C1(net938),
    .X(_00099_));
 sky130_fd_sc_hd__a21boi_1 _17427_ (.A1(net27),
    .A2(net28),
    .B1_N(net222),
    .Y(_08562_));
 sky130_fd_sc_hd__and4_4 _17428_ (.A(net67),
    .B(net933),
    .C(_08390_),
    .D(_08562_),
    .X(_00100_));
 sky130_fd_sc_hd__or3_4 _17429_ (.A(net69),
    .B(_08393_),
    .C(net265),
    .X(_08563_));
 sky130_fd_sc_hd__mux2_1 _17430_ (.A0(net35),
    .A1(\op_code[0] ),
    .S(_08563_),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _17431_ (.A0(net46),
    .A1(\op_code[1] ),
    .S(_08563_),
    .X(_00102_));
 sky130_fd_sc_hd__mux2_1 _17432_ (.A0(net57),
    .A1(net316),
    .S(_08563_),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_1 _17433_ (.A0(net60),
    .A1(net315),
    .S(_08563_),
    .X(_00104_));
 sky130_fd_sc_hd__dfxtp_2 _17434_ (.CLK(clknet_4_0_0_clk),
    .D(_00004_),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_4 _17435_ (.CLK(clknet_4_8_0_clk),
    .D(_00005_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_4 _17436_ (.CLK(clknet_4_8_0_clk),
    .D(_00006_),
    .Q(net105));
 sky130_fd_sc_hd__dfxtp_4 _17437_ (.CLK(clknet_4_14_0_clk),
    .D(_00007_),
    .Q(net108));
 sky130_fd_sc_hd__dfxtp_4 _17438_ (.CLK(clknet_4_9_0_clk),
    .D(_00008_),
    .Q(net109));
 sky130_fd_sc_hd__dfxtp_2 _17439_ (.CLK(clknet_4_0_0_clk),
    .D(_00009_),
    .Q(net110));
 sky130_fd_sc_hd__dfxtp_4 _17440_ (.CLK(clknet_4_2_0_clk),
    .D(_00010_),
    .Q(net111));
 sky130_fd_sc_hd__dfxtp_4 _17441_ (.CLK(clknet_4_2_0_clk),
    .D(_00011_),
    .Q(net112));
 sky130_fd_sc_hd__dfxtp_4 _17442_ (.CLK(clknet_4_9_0_clk),
    .D(_00012_),
    .Q(net113));
 sky130_fd_sc_hd__dfxtp_4 _17443_ (.CLK(clknet_4_9_0_clk),
    .D(_00013_),
    .Q(net114));
 sky130_fd_sc_hd__dfxtp_4 _17444_ (.CLK(clknet_4_13_0_clk),
    .D(_00014_),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_2 _17445_ (.CLK(clknet_4_4_0_clk),
    .D(_00015_),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_4 _17446_ (.CLK(clknet_4_1_0_clk),
    .D(_00016_),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_4 _17447_ (.CLK(clknet_4_2_0_clk),
    .D(_00017_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_2 _17448_ (.CLK(clknet_4_1_0_clk),
    .D(_00018_),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_4 _17449_ (.CLK(clknet_4_1_0_clk),
    .D(_00019_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_2 _17450_ (.CLK(clknet_4_4_0_clk),
    .D(_00020_),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_2 _17451_ (.CLK(clknet_4_4_0_clk),
    .D(_00021_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_2 _17452_ (.CLK(clknet_4_5_0_clk),
    .D(_00022_),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_2 _17453_ (.CLK(clknet_4_5_0_clk),
    .D(_00023_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_2 _17454_ (.CLK(clknet_4_4_0_clk),
    .D(_00024_),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_2 _17455_ (.CLK(clknet_4_5_0_clk),
    .D(_00025_),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_2 _17456_ (.CLK(clknet_4_5_0_clk),
    .D(_00026_),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_4 _17457_ (.CLK(clknet_4_7_0_clk),
    .D(_00027_),
    .Q(net98));
 sky130_fd_sc_hd__dfxtp_2 _17458_ (.CLK(clknet_4_4_0_clk),
    .D(_00028_),
    .Q(net99));
 sky130_fd_sc_hd__dfxtp_4 _17459_ (.CLK(clknet_4_7_0_clk),
    .D(_00029_),
    .Q(net100));
 sky130_fd_sc_hd__dfxtp_4 _17460_ (.CLK(clknet_4_4_0_clk),
    .D(_00030_),
    .Q(net101));
 sky130_fd_sc_hd__dfxtp_4 _17461_ (.CLK(clknet_4_6_0_clk),
    .D(_00031_),
    .Q(net102));
 sky130_fd_sc_hd__dfxtp_4 _17462_ (.CLK(clknet_4_4_0_clk),
    .D(_00032_),
    .Q(net103));
 sky130_fd_sc_hd__dfxtp_4 _17463_ (.CLK(clknet_4_6_0_clk),
    .D(_00033_),
    .Q(net104));
 sky130_fd_sc_hd__dfxtp_4 _17464_ (.CLK(clknet_4_1_0_clk),
    .D(_00034_),
    .Q(net106));
 sky130_fd_sc_hd__dfxtp_4 _17465_ (.CLK(clknet_4_7_0_clk),
    .D(_00035_),
    .Q(net107));
 sky130_fd_sc_hd__dfxtp_2 _17466_ (.CLK(clknet_4_10_0_clk),
    .D(net914),
    .Q(net70));
 sky130_fd_sc_hd__dfxtp_4 _17467_ (.CLK(clknet_4_10_0_clk),
    .D(net906),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_2 _17468_ (.CLK(clknet_4_10_0_clk),
    .D(net899),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_4 _17469_ (.CLK(clknet_4_10_0_clk),
    .D(net889),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_4 _17470_ (.CLK(clknet_4_11_0_clk),
    .D(\salida[0] ),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_4 _17471_ (.CLK(clknet_4_10_0_clk),
    .D(\salida[1] ),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_4 _17472_ (.CLK(clknet_4_10_0_clk),
    .D(\salida[2] ),
    .Q(net78));
 sky130_fd_sc_hd__dfxtp_4 _17473_ (.CLK(clknet_4_10_0_clk),
    .D(\salida[3] ),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_4 _17474_ (.CLK(clknet_4_11_0_clk),
    .D(\op_code[0] ),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_4 _17475_ (.CLK(clknet_4_11_0_clk),
    .D(\op_code[1] ),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_4 _17476_ (.CLK(clknet_4_11_0_clk),
    .D(\op_code[2] ),
    .Q(net71));
 sky130_fd_sc_hd__dfxtp_4 _17477_ (.CLK(clknet_4_11_0_clk),
    .D(net315),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_4 _17478_ (.CLK(clknet_4_14_0_clk),
    .D(_00036_),
    .Q(\ApproximateM_inst.lob_16.lob1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_4 _17479_ (.CLK(clknet_4_14_0_clk),
    .D(_00037_),
    .Q(\ApproximateM_inst.lob_16.lob1.genblk1[1].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_4 _17480_ (.CLK(clknet_4_12_0_clk),
    .D(_00038_),
    .Q(\ApproximateM_inst.lob_16.lob1.genblk1[2].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_1 _17481_ (.CLK(clknet_4_12_0_clk),
    .D(_00039_),
    .Q(\ApproximateM_inst.lob_16.lob1.genblk1[3].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_1 _17482_ (.CLK(clknet_4_14_0_clk),
    .D(_00040_),
    .Q(\ApproximateM_inst.lob_16.lob1.genblk1[4].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_1 _17483_ (.CLK(clknet_4_15_0_clk),
    .D(_00041_),
    .Q(\ApproximateM_inst.lob_16.lob1.genblk1[5].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_4 _17484_ (.CLK(clknet_4_15_0_clk),
    .D(_00042_),
    .Q(\ApproximateM_inst.lob_16.lob1.genblk1[6].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_4 _17485_ (.CLK(clknet_4_14_0_clk),
    .D(_00043_),
    .Q(\ApproximateM_inst.lob_16.lob1.genblk1[7].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_1 _17486_ (.CLK(clknet_4_15_0_clk),
    .D(_00044_),
    .Q(\ApproximateM_inst.lob_16.lob1.genblk1[8].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_4 _17487_ (.CLK(clknet_4_12_0_clk),
    .D(_00045_),
    .Q(\ApproximateM_inst.lob_16.lob1.genblk1[9].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_4 _17488_ (.CLK(clknet_4_15_0_clk),
    .D(_00046_),
    .Q(\ApproximateM_inst.lob_16.lob1.genblk1[10].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_1 _17489_ (.CLK(clknet_4_15_0_clk),
    .D(_00047_),
    .Q(\ApproximateM_inst.lob_16.lob1.genblk1[11].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_1 _17490_ (.CLK(clknet_4_15_0_clk),
    .D(_00048_),
    .Q(\ApproximateM_inst.lob_16.lob1.genblk1[12].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_1 _17491_ (.CLK(clknet_4_15_0_clk),
    .D(_00049_),
    .Q(\ApproximateM_inst.lob_16.lob1.genblk1[13].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_4 _17492_ (.CLK(clknet_4_15_0_clk),
    .D(_00050_),
    .Q(\ApproximateM_inst.lob_16.lob1.genblk1[14].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_4 _17493_ (.CLK(clknet_4_14_0_clk),
    .D(_00051_),
    .Q(\ApproximateM_inst.lob_16.lob1.genblk2.mux_final.sel ));
 sky130_fd_sc_hd__dfxtp_1 _17494_ (.CLK(clknet_4_15_0_clk),
    .D(_00052_),
    .Q(\cla_inst.in1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _17495_ (.CLK(clknet_4_14_0_clk),
    .D(_00053_),
    .Q(\cla_inst.in1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _17496_ (.CLK(clknet_4_15_0_clk),
    .D(_00054_),
    .Q(\cla_inst.in1[18] ));
 sky130_fd_sc_hd__dfxtp_2 _17497_ (.CLK(clknet_4_12_0_clk),
    .D(_00055_),
    .Q(\cla_inst.in1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _17498_ (.CLK(clknet_4_12_0_clk),
    .D(_00056_),
    .Q(\cla_inst.in1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _17499_ (.CLK(clknet_4_12_0_clk),
    .D(_00057_),
    .Q(\cla_inst.in1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _17500_ (.CLK(clknet_4_12_0_clk),
    .D(_00058_),
    .Q(\cla_inst.in1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _17501_ (.CLK(clknet_4_13_0_clk),
    .D(_00059_),
    .Q(\cla_inst.in1[23] ));
 sky130_fd_sc_hd__dfxtp_2 _17502_ (.CLK(clknet_4_12_0_clk),
    .D(_00060_),
    .Q(\cla_inst.in1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _17503_ (.CLK(clknet_4_13_0_clk),
    .D(_00061_),
    .Q(\cla_inst.in1[25] ));
 sky130_fd_sc_hd__dfxtp_4 _17504_ (.CLK(clknet_4_13_0_clk),
    .D(_00062_),
    .Q(\cla_inst.in1[26] ));
 sky130_fd_sc_hd__dfxtp_4 _17505_ (.CLK(clknet_4_13_0_clk),
    .D(_00063_),
    .Q(\cla_inst.in1[27] ));
 sky130_fd_sc_hd__dfxtp_4 _17506_ (.CLK(clknet_4_13_0_clk),
    .D(_00064_),
    .Q(\cla_inst.in1[28] ));
 sky130_fd_sc_hd__dfxtp_4 _17507_ (.CLK(clknet_4_13_0_clk),
    .D(_00065_),
    .Q(\cla_inst.in1[29] ));
 sky130_fd_sc_hd__dfxtp_2 _17508_ (.CLK(clknet_4_13_0_clk),
    .D(_00066_),
    .Q(\cla_inst.in1[30] ));
 sky130_fd_sc_hd__dfxtp_2 _17509_ (.CLK(clknet_4_13_0_clk),
    .D(_00067_),
    .Q(\cla_inst.in1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _17510_ (.CLK(clknet_4_8_0_clk),
    .D(_00068_),
    .Q(\ApproximateM_inst.lob_16.lob2.mux.sel ));
 sky130_fd_sc_hd__dfxtp_4 _17511_ (.CLK(clknet_4_14_0_clk),
    .D(_00069_),
    .Q(\ApproximateM_inst.lob_16.lob2.genblk1[1].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_1 _17512_ (.CLK(clknet_4_8_0_clk),
    .D(_00070_),
    .Q(\ApproximateM_inst.lob_16.lob2.genblk1[2].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_1 _17513_ (.CLK(clknet_4_8_0_clk),
    .D(_00071_),
    .Q(\ApproximateM_inst.lob_16.lob2.genblk1[3].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_1 _17514_ (.CLK(clknet_4_14_0_clk),
    .D(_00072_),
    .Q(\ApproximateM_inst.lob_16.lob2.genblk1[4].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_1 _17515_ (.CLK(clknet_4_15_0_clk),
    .D(_00073_),
    .Q(\ApproximateM_inst.lob_16.lob2.genblk1[5].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_4 _17516_ (.CLK(clknet_4_15_0_clk),
    .D(_00074_),
    .Q(\ApproximateM_inst.lob_16.lob2.genblk1[6].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_4 _17517_ (.CLK(clknet_4_8_0_clk),
    .D(_00075_),
    .Q(\ApproximateM_inst.lob_16.lob2.genblk1[7].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_1 _17518_ (.CLK(clknet_4_12_0_clk),
    .D(_00076_),
    .Q(\ApproximateM_inst.lob_16.lob2.genblk1[8].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_4 _17519_ (.CLK(clknet_4_12_0_clk),
    .D(_00077_),
    .Q(\ApproximateM_inst.lob_16.lob2.genblk1[9].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_4 _17520_ (.CLK(clknet_4_15_0_clk),
    .D(_00078_),
    .Q(\ApproximateM_inst.lob_16.lob2.genblk1[10].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_4 _17521_ (.CLK(clknet_4_15_0_clk),
    .D(_00079_),
    .Q(\ApproximateM_inst.lob_16.lob2.genblk1[11].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_1 _17522_ (.CLK(clknet_4_15_0_clk),
    .D(_00080_),
    .Q(\ApproximateM_inst.lob_16.lob2.genblk1[12].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_1 _17523_ (.CLK(clknet_4_15_0_clk),
    .D(_00081_),
    .Q(\ApproximateM_inst.lob_16.lob2.genblk1[13].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_1 _17524_ (.CLK(clknet_4_15_0_clk),
    .D(_00082_),
    .Q(\ApproximateM_inst.lob_16.lob2.genblk1[14].genblk1.mux.sel ));
 sky130_fd_sc_hd__dfxtp_2 _17525_ (.CLK(clknet_4_15_0_clk),
    .D(_00083_),
    .Q(\ApproximateM_inst.lob_16.lob2.genblk2.mux_final.sel ));
 sky130_fd_sc_hd__dfxtp_1 _17526_ (.CLK(clknet_4_15_0_clk),
    .D(_00084_),
    .Q(\cla_inst.in2[16] ));
 sky130_fd_sc_hd__dfxtp_1 _17527_ (.CLK(clknet_4_15_0_clk),
    .D(_00085_),
    .Q(\cla_inst.in2[17] ));
 sky130_fd_sc_hd__dfxtp_4 _17528_ (.CLK(clknet_4_14_0_clk),
    .D(_00086_),
    .Q(\cla_inst.in2[18] ));
 sky130_fd_sc_hd__dfxtp_1 _17529_ (.CLK(clknet_4_15_0_clk),
    .D(_00087_),
    .Q(\cla_inst.in2[19] ));
 sky130_fd_sc_hd__dfxtp_4 _17530_ (.CLK(clknet_4_12_0_clk),
    .D(_00088_),
    .Q(\cla_inst.in2[20] ));
 sky130_fd_sc_hd__dfxtp_4 _17531_ (.CLK(clknet_4_12_0_clk),
    .D(_00089_),
    .Q(\cla_inst.in2[21] ));
 sky130_fd_sc_hd__dfxtp_4 _17532_ (.CLK(clknet_4_12_0_clk),
    .D(_00090_),
    .Q(\cla_inst.in2[22] ));
 sky130_fd_sc_hd__dfxtp_4 _17533_ (.CLK(clknet_4_12_0_clk),
    .D(_00091_),
    .Q(\cla_inst.in2[23] ));
 sky130_fd_sc_hd__dfxtp_1 _17534_ (.CLK(clknet_4_13_0_clk),
    .D(_00092_),
    .Q(\cla_inst.in2[24] ));
 sky130_fd_sc_hd__dfxtp_1 _17535_ (.CLK(clknet_4_13_0_clk),
    .D(_00093_),
    .Q(\cla_inst.in2[25] ));
 sky130_fd_sc_hd__dfxtp_1 _17536_ (.CLK(clknet_4_13_0_clk),
    .D(_00094_),
    .Q(\cla_inst.in2[26] ));
 sky130_fd_sc_hd__dfxtp_1 _17537_ (.CLK(clknet_4_13_0_clk),
    .D(_00095_),
    .Q(\cla_inst.in2[27] ));
 sky130_fd_sc_hd__dfxtp_2 _17538_ (.CLK(clknet_4_13_0_clk),
    .D(_00096_),
    .Q(\cla_inst.in2[28] ));
 sky130_fd_sc_hd__dfxtp_4 _17539_ (.CLK(clknet_4_0_0_clk),
    .D(_00097_),
    .Q(\cla_inst.in2[29] ));
 sky130_fd_sc_hd__dfxtp_2 _17540_ (.CLK(clknet_4_0_0_clk),
    .D(_00098_),
    .Q(\cla_inst.in2[30] ));
 sky130_fd_sc_hd__dfxtp_1 _17541_ (.CLK(clknet_4_0_0_clk),
    .D(_00099_),
    .Q(\cla_inst.in2[31] ));
 sky130_fd_sc_hd__dfxtp_1 _17542_ (.CLK(clknet_4_3_0_clk),
    .D(_00100_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_2 _17543_ (.CLK(clknet_4_11_0_clk),
    .D(_08684_),
    .Q(\salida[0] ));
 sky130_fd_sc_hd__dfxtp_2 _17544_ (.CLK(clknet_4_10_0_clk),
    .D(_08695_),
    .Q(\salida[1] ));
 sky130_fd_sc_hd__dfxtp_2 _17545_ (.CLK(clknet_4_10_0_clk),
    .D(_08706_),
    .Q(\salida[2] ));
 sky130_fd_sc_hd__dfxtp_4 _17546_ (.CLK(clknet_4_10_0_clk),
    .D(_08709_),
    .Q(\salida[3] ));
 sky130_fd_sc_hd__dfxtp_1 _17547_ (.CLK(clknet_4_9_0_clk),
    .D(_08710_),
    .Q(\salida[4] ));
 sky130_fd_sc_hd__dfxtp_1 _17548_ (.CLK(clknet_4_2_0_clk),
    .D(_08711_),
    .Q(\salida[5] ));
 sky130_fd_sc_hd__dfxtp_1 _17549_ (.CLK(clknet_4_2_0_clk),
    .D(_08712_),
    .Q(\salida[6] ));
 sky130_fd_sc_hd__dfxtp_1 _17550_ (.CLK(clknet_4_9_0_clk),
    .D(_08713_),
    .Q(\salida[7] ));
 sky130_fd_sc_hd__dfxtp_1 _17551_ (.CLK(clknet_4_10_0_clk),
    .D(_08714_),
    .Q(\salida[8] ));
 sky130_fd_sc_hd__dfxtp_1 _17552_ (.CLK(clknet_4_8_0_clk),
    .D(_08715_),
    .Q(\salida[9] ));
 sky130_fd_sc_hd__dfxtp_1 _17553_ (.CLK(clknet_4_11_0_clk),
    .D(_08685_),
    .Q(\salida[10] ));
 sky130_fd_sc_hd__dfxtp_2 _17554_ (.CLK(clknet_4_11_0_clk),
    .D(_08686_),
    .Q(\salida[11] ));
 sky130_fd_sc_hd__dfxtp_1 _17555_ (.CLK(clknet_4_3_0_clk),
    .D(_08687_),
    .Q(\salida[12] ));
 sky130_fd_sc_hd__dfxtp_1 _17556_ (.CLK(clknet_4_2_0_clk),
    .D(_08688_),
    .Q(\salida[13] ));
 sky130_fd_sc_hd__dfxtp_1 _17557_ (.CLK(clknet_4_0_0_clk),
    .D(_08689_),
    .Q(\salida[14] ));
 sky130_fd_sc_hd__dfxtp_1 _17558_ (.CLK(clknet_4_2_0_clk),
    .D(_08690_),
    .Q(\salida[15] ));
 sky130_fd_sc_hd__dfxtp_1 _17559_ (.CLK(clknet_4_4_0_clk),
    .D(_08691_),
    .Q(\salida[16] ));
 sky130_fd_sc_hd__dfxtp_1 _17560_ (.CLK(clknet_4_6_0_clk),
    .D(_08692_),
    .Q(\salida[17] ));
 sky130_fd_sc_hd__dfxtp_1 _17561_ (.CLK(clknet_4_4_0_clk),
    .D(_08693_),
    .Q(\salida[18] ));
 sky130_fd_sc_hd__dfxtp_1 _17562_ (.CLK(clknet_4_7_0_clk),
    .D(_08694_),
    .Q(\salida[19] ));
 sky130_fd_sc_hd__dfxtp_1 _17563_ (.CLK(clknet_4_5_0_clk),
    .D(_08696_),
    .Q(\salida[20] ));
 sky130_fd_sc_hd__dfxtp_1 _17564_ (.CLK(clknet_4_5_0_clk),
    .D(_08697_),
    .Q(\salida[21] ));
 sky130_fd_sc_hd__dfxtp_1 _17565_ (.CLK(clknet_4_5_0_clk),
    .D(_08698_),
    .Q(\salida[22] ));
 sky130_fd_sc_hd__dfxtp_1 _17566_ (.CLK(clknet_4_7_0_clk),
    .D(_08699_),
    .Q(\salida[23] ));
 sky130_fd_sc_hd__dfxtp_1 _17567_ (.CLK(clknet_4_5_0_clk),
    .D(_08700_),
    .Q(\salida[24] ));
 sky130_fd_sc_hd__dfxtp_1 _17568_ (.CLK(clknet_4_4_0_clk),
    .D(_08701_),
    .Q(\salida[25] ));
 sky130_fd_sc_hd__dfxtp_1 _17569_ (.CLK(clknet_4_6_0_clk),
    .D(_08702_),
    .Q(\salida[26] ));
 sky130_fd_sc_hd__dfxtp_1 _17570_ (.CLK(clknet_4_6_0_clk),
    .D(_08703_),
    .Q(\salida[27] ));
 sky130_fd_sc_hd__dfxtp_1 _17571_ (.CLK(clknet_4_6_0_clk),
    .D(_08704_),
    .Q(\salida[28] ));
 sky130_fd_sc_hd__dfxtp_1 _17572_ (.CLK(clknet_4_3_0_clk),
    .D(_08705_),
    .Q(\salida[29] ));
 sky130_fd_sc_hd__dfxtp_1 _17573_ (.CLK(clknet_4_3_0_clk),
    .D(_08707_),
    .Q(\salida[30] ));
 sky130_fd_sc_hd__dfxtp_1 _17574_ (.CLK(clknet_4_3_0_clk),
    .D(_08708_),
    .Q(\salida[31] ));
 sky130_fd_sc_hd__dfxtp_1 _17575_ (.CLK(clknet_4_13_0_clk),
    .D(_08716_),
    .Q(\salida[32] ));
 sky130_fd_sc_hd__dfxtp_1 _17576_ (.CLK(clknet_4_8_0_clk),
    .D(_08653_),
    .Q(\salida[33] ));
 sky130_fd_sc_hd__dfxtp_1 _17577_ (.CLK(clknet_4_14_0_clk),
    .D(_08664_),
    .Q(\salida[34] ));
 sky130_fd_sc_hd__dfxtp_1 _17578_ (.CLK(clknet_4_14_0_clk),
    .D(_08675_),
    .Q(\salida[35] ));
 sky130_fd_sc_hd__dfxtp_1 _17579_ (.CLK(clknet_4_8_0_clk),
    .D(_08677_),
    .Q(\salida[36] ));
 sky130_fd_sc_hd__dfxtp_1 _17580_ (.CLK(clknet_4_0_0_clk),
    .D(_08678_),
    .Q(\salida[37] ));
 sky130_fd_sc_hd__dfxtp_1 _17581_ (.CLK(clknet_4_14_0_clk),
    .D(_08679_),
    .Q(\salida[38] ));
 sky130_fd_sc_hd__dfxtp_1 _17582_ (.CLK(clknet_4_8_0_clk),
    .D(_08680_),
    .Q(\salida[39] ));
 sky130_fd_sc_hd__dfxtp_1 _17583_ (.CLK(clknet_4_14_0_clk),
    .D(_08681_),
    .Q(\salida[40] ));
 sky130_fd_sc_hd__dfxtp_1 _17584_ (.CLK(clknet_4_8_0_clk),
    .D(_08682_),
    .Q(\salida[41] ));
 sky130_fd_sc_hd__dfxtp_1 _17585_ (.CLK(clknet_4_9_0_clk),
    .D(_08683_),
    .Q(\salida[42] ));
 sky130_fd_sc_hd__dfxtp_1 _17586_ (.CLK(clknet_4_1_0_clk),
    .D(_08654_),
    .Q(\salida[43] ));
 sky130_fd_sc_hd__dfxtp_1 _17587_ (.CLK(clknet_4_1_0_clk),
    .D(_08655_),
    .Q(\salida[44] ));
 sky130_fd_sc_hd__dfxtp_1 _17588_ (.CLK(clknet_4_0_0_clk),
    .D(_08656_),
    .Q(\salida[45] ));
 sky130_fd_sc_hd__dfxtp_1 _17589_ (.CLK(clknet_4_1_0_clk),
    .D(_08657_),
    .Q(\salida[46] ));
 sky130_fd_sc_hd__dfxtp_1 _17590_ (.CLK(clknet_4_1_0_clk),
    .D(_08658_),
    .Q(\salida[47] ));
 sky130_fd_sc_hd__dfxtp_1 _17591_ (.CLK(clknet_4_4_0_clk),
    .D(_08659_),
    .Q(\salida[48] ));
 sky130_fd_sc_hd__dfxtp_1 _17592_ (.CLK(clknet_4_4_0_clk),
    .D(_08660_),
    .Q(\salida[49] ));
 sky130_fd_sc_hd__dfxtp_1 _17593_ (.CLK(clknet_4_5_0_clk),
    .D(_08661_),
    .Q(\salida[50] ));
 sky130_fd_sc_hd__dfxtp_1 _17594_ (.CLK(clknet_4_5_0_clk),
    .D(_08662_),
    .Q(\salida[51] ));
 sky130_fd_sc_hd__dfxtp_1 _17595_ (.CLK(clknet_4_4_0_clk),
    .D(_08663_),
    .Q(\salida[52] ));
 sky130_fd_sc_hd__dfxtp_1 _17596_ (.CLK(clknet_4_5_0_clk),
    .D(_08665_),
    .Q(\salida[53] ));
 sky130_fd_sc_hd__dfxtp_1 _17597_ (.CLK(clknet_4_7_0_clk),
    .D(_08666_),
    .Q(\salida[54] ));
 sky130_fd_sc_hd__dfxtp_1 _17598_ (.CLK(clknet_4_7_0_clk),
    .D(_08667_),
    .Q(\salida[55] ));
 sky130_fd_sc_hd__dfxtp_1 _17599_ (.CLK(clknet_4_4_0_clk),
    .D(_08668_),
    .Q(\salida[56] ));
 sky130_fd_sc_hd__dfxtp_1 _17600_ (.CLK(clknet_4_6_0_clk),
    .D(_08669_),
    .Q(\salida[57] ));
 sky130_fd_sc_hd__dfxtp_1 _17601_ (.CLK(clknet_4_6_0_clk),
    .D(_08670_),
    .Q(\salida[58] ));
 sky130_fd_sc_hd__dfxtp_1 _17602_ (.CLK(clknet_4_6_0_clk),
    .D(_08671_),
    .Q(\salida[59] ));
 sky130_fd_sc_hd__dfxtp_1 _17603_ (.CLK(clknet_4_4_0_clk),
    .D(_08672_),
    .Q(\salida[60] ));
 sky130_fd_sc_hd__dfxtp_1 _17604_ (.CLK(clknet_4_6_0_clk),
    .D(_08673_),
    .Q(\salida[61] ));
 sky130_fd_sc_hd__dfxtp_1 _17605_ (.CLK(clknet_4_1_0_clk),
    .D(_08674_),
    .Q(\salida[62] ));
 sky130_fd_sc_hd__dfxtp_1 _17606_ (.CLK(clknet_4_1_0_clk),
    .D(_08676_),
    .Q(\salida[63] ));
 sky130_fd_sc_hd__dfxtp_4 _17607_ (.CLK(clknet_4_9_0_clk),
    .D(_00101_),
    .Q(\op_code[0] ));
 sky130_fd_sc_hd__dfxtp_4 _17608_ (.CLK(clknet_4_9_0_clk),
    .D(_00102_),
    .Q(\op_code[1] ));
 sky130_fd_sc_hd__dfxtp_4 _17609_ (.CLK(clknet_4_9_0_clk),
    .D(_00103_),
    .Q(\op_code[2] ));
 sky130_fd_sc_hd__dfxtp_2 _17610_ (.CLK(clknet_4_9_0_clk),
    .D(_00104_),
    .Q(\op_code[3] ));
 sky130_fd_sc_hd__dfxtp_1 _17611_ (.CLK(clknet_4_11_0_clk),
    .D(_00000_),
    .Q(\sel_op[0] ));
 sky130_fd_sc_hd__dfxtp_1 _17612_ (.CLK(clknet_4_11_0_clk),
    .D(_00001_),
    .Q(\sel_op[1] ));
 sky130_fd_sc_hd__dfxtp_2 _17613_ (.CLK(clknet_4_11_0_clk),
    .D(_00002_),
    .Q(\sel_op[2] ));
 sky130_fd_sc_hd__dfxtp_4 _17614_ (.CLK(clknet_4_11_0_clk),
    .D(_00003_),
    .Q(\sel_op[3] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__buf_4 fanout123 (.A(net126),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_4 fanout124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__buf_4 fanout125 (.A(net126),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_4 fanout126 (.A(_08406_),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_8 fanout127 (.A(net130),
    .X(net127));
 sky130_fd_sc_hd__buf_4 fanout128 (.A(net129),
    .X(net128));
 sky130_fd_sc_hd__buf_4 fanout129 (.A(net130),
    .X(net129));
 sky130_fd_sc_hd__buf_4 fanout130 (.A(_08394_),
    .X(net130));
 sky130_fd_sc_hd__buf_8 fanout131 (.A(net132),
    .X(net131));
 sky130_fd_sc_hd__buf_6 fanout132 (.A(_06447_),
    .X(net132));
 sky130_fd_sc_hd__buf_6 fanout133 (.A(net135),
    .X(net133));
 sky130_fd_sc_hd__buf_6 fanout134 (.A(net135),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_16 fanout135 (.A(_06386_),
    .X(net135));
 sky130_fd_sc_hd__buf_12 fanout136 (.A(_06234_),
    .X(net136));
 sky130_fd_sc_hd__buf_4 fanout137 (.A(_06234_),
    .X(net137));
 sky130_fd_sc_hd__buf_6 fanout138 (.A(_06104_),
    .X(net138));
 sky130_fd_sc_hd__buf_12 fanout140 (.A(_06097_),
    .X(net140));
 sky130_fd_sc_hd__buf_8 fanout141 (.A(net142),
    .X(net141));
 sky130_fd_sc_hd__buf_12 fanout142 (.A(_06047_),
    .X(net142));
 sky130_fd_sc_hd__buf_4 fanout143 (.A(net144),
    .X(net143));
 sky130_fd_sc_hd__buf_6 fanout144 (.A(_06041_),
    .X(net144));
 sky130_fd_sc_hd__buf_6 fanout145 (.A(net147),
    .X(net145));
 sky130_fd_sc_hd__buf_4 fanout146 (.A(net147),
    .X(net146));
 sky130_fd_sc_hd__buf_6 fanout147 (.A(_05990_),
    .X(net147));
 sky130_fd_sc_hd__buf_4 fanout148 (.A(_05985_),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_2 fanout149 (.A(_05985_),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_4 fanout150 (.A(_05924_),
    .X(net150));
 sky130_fd_sc_hd__buf_4 fanout151 (.A(_05923_),
    .X(net151));
 sky130_fd_sc_hd__buf_4 fanout152 (.A(_05923_),
    .X(net152));
 sky130_fd_sc_hd__buf_8 fanout153 (.A(_05919_),
    .X(net153));
 sky130_fd_sc_hd__buf_6 fanout154 (.A(net155),
    .X(net154));
 sky130_fd_sc_hd__buf_6 fanout155 (.A(_05900_),
    .X(net155));
 sky130_fd_sc_hd__buf_4 fanout156 (.A(net159),
    .X(net156));
 sky130_fd_sc_hd__buf_2 fanout157 (.A(net159),
    .X(net157));
 sky130_fd_sc_hd__buf_4 fanout158 (.A(net159),
    .X(net158));
 sky130_fd_sc_hd__buf_2 fanout159 (.A(_08523_),
    .X(net159));
 sky130_fd_sc_hd__buf_4 fanout160 (.A(_08523_),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_4 fanout161 (.A(net163),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_2 fanout162 (.A(net163),
    .X(net162));
 sky130_fd_sc_hd__buf_4 fanout163 (.A(_08522_),
    .X(net163));
 sky130_fd_sc_hd__buf_4 fanout164 (.A(_08482_),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_4 fanout165 (.A(_08482_),
    .X(net165));
 sky130_fd_sc_hd__buf_4 fanout166 (.A(_08482_),
    .X(net166));
 sky130_fd_sc_hd__buf_2 fanout167 (.A(_08482_),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_4 fanout168 (.A(_07129_),
    .X(net168));
 sky130_fd_sc_hd__buf_4 fanout169 (.A(_06907_),
    .X(net169));
 sky130_fd_sc_hd__buf_4 fanout170 (.A(_06906_),
    .X(net170));
 sky130_fd_sc_hd__buf_4 fanout171 (.A(_06806_),
    .X(net171));
 sky130_fd_sc_hd__buf_6 fanout172 (.A(_06805_),
    .X(net172));
 sky130_fd_sc_hd__buf_6 fanout173 (.A(net174),
    .X(net173));
 sky130_fd_sc_hd__buf_6 fanout174 (.A(_06732_),
    .X(net174));
 sky130_fd_sc_hd__buf_4 fanout175 (.A(net176),
    .X(net175));
 sky130_fd_sc_hd__buf_4 fanout176 (.A(_06644_),
    .X(net176));
 sky130_fd_sc_hd__buf_6 fanout177 (.A(_06643_),
    .X(net177));
 sky130_fd_sc_hd__buf_4 fanout178 (.A(_06643_),
    .X(net178));
 sky130_fd_sc_hd__buf_4 fanout179 (.A(net181),
    .X(net179));
 sky130_fd_sc_hd__buf_2 fanout180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_4 fanout181 (.A(_06618_),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_8 fanout182 (.A(_06617_),
    .X(net182));
 sky130_fd_sc_hd__buf_6 fanout183 (.A(_06553_),
    .X(net183));
 sky130_fd_sc_hd__buf_8 fanout184 (.A(_06552_),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_8 fanout185 (.A(_06531_),
    .X(net185));
 sky130_fd_sc_hd__buf_4 fanout186 (.A(_06531_),
    .X(net186));
 sky130_fd_sc_hd__buf_4 fanout187 (.A(_06465_),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_16 fanout188 (.A(_06464_),
    .X(net188));
 sky130_fd_sc_hd__buf_8 fanout189 (.A(net190),
    .X(net189));
 sky130_fd_sc_hd__buf_6 fanout190 (.A(_06373_),
    .X(net190));
 sky130_fd_sc_hd__buf_8 fanout191 (.A(net192),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_8 fanout192 (.A(_06314_),
    .X(net192));
 sky130_fd_sc_hd__buf_6 fanout194 (.A(_06304_),
    .X(net194));
 sky130_fd_sc_hd__buf_2 fanout195 (.A(_06304_),
    .X(net195));
 sky130_fd_sc_hd__buf_6 fanout196 (.A(_06247_),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_16 fanout198 (.A(_06183_),
    .X(net198));
 sky130_fd_sc_hd__buf_4 fanout199 (.A(_06183_),
    .X(net199));
 sky130_fd_sc_hd__buf_12 fanout200 (.A(_06176_),
    .X(net200));
 sky130_fd_sc_hd__buf_4 fanout201 (.A(_06176_),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_8 fanout202 (.A(net203),
    .X(net202));
 sky130_fd_sc_hd__buf_6 fanout203 (.A(_05939_),
    .X(net203));
 sky130_fd_sc_hd__buf_4 fanout204 (.A(_04528_),
    .X(net204));
 sky130_fd_sc_hd__buf_4 fanout205 (.A(_03686_),
    .X(net205));
 sky130_fd_sc_hd__buf_6 fanout206 (.A(net207),
    .X(net206));
 sky130_fd_sc_hd__buf_6 fanout207 (.A(_02648_),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_8 fanout208 (.A(net209),
    .X(net208));
 sky130_fd_sc_hd__buf_6 fanout209 (.A(_02644_),
    .X(net209));
 sky130_fd_sc_hd__buf_4 fanout210 (.A(_02644_),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_4 fanout211 (.A(_02644_),
    .X(net211));
 sky130_fd_sc_hd__buf_4 fanout212 (.A(net215),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_4 fanout213 (.A(net215),
    .X(net213));
 sky130_fd_sc_hd__buf_6 fanout214 (.A(net215),
    .X(net214));
 sky130_fd_sc_hd__buf_4 fanout215 (.A(net216),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_4 fanout218 (.A(_08404_),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_4 fanout219 (.A(_08404_),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_4 fanout220 (.A(_08404_),
    .X(net220));
 sky130_fd_sc_hd__buf_2 fanout221 (.A(_08404_),
    .X(net221));
 sky130_fd_sc_hd__buf_4 fanout223 (.A(net224),
    .X(net223));
 sky130_fd_sc_hd__buf_6 fanout224 (.A(_06711_),
    .X(net224));
 sky130_fd_sc_hd__buf_12 fanout225 (.A(net226),
    .X(net225));
 sky130_fd_sc_hd__buf_4 fanout226 (.A(net227),
    .X(net226));
 sky130_fd_sc_hd__buf_4 fanout227 (.A(_06179_),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_8 fanout228 (.A(net229),
    .X(net228));
 sky130_fd_sc_hd__buf_6 fanout229 (.A(_05952_),
    .X(net229));
 sky130_fd_sc_hd__buf_6 fanout230 (.A(_05951_),
    .X(net230));
 sky130_fd_sc_hd__buf_4 fanout231 (.A(net234),
    .X(net231));
 sky130_fd_sc_hd__buf_4 fanout232 (.A(net233),
    .X(net232));
 sky130_fd_sc_hd__buf_4 fanout233 (.A(net234),
    .X(net233));
 sky130_fd_sc_hd__buf_4 fanout234 (.A(_05947_),
    .X(net234));
 sky130_fd_sc_hd__buf_6 fanout235 (.A(_05945_),
    .X(net235));
 sky130_fd_sc_hd__buf_4 fanout236 (.A(net237),
    .X(net236));
 sky130_fd_sc_hd__buf_6 fanout237 (.A(_05944_),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_8 fanout238 (.A(net239),
    .X(net238));
 sky130_fd_sc_hd__buf_4 fanout239 (.A(net240),
    .X(net239));
 sky130_fd_sc_hd__buf_6 fanout240 (.A(_05941_),
    .X(net240));
 sky130_fd_sc_hd__buf_6 fanout241 (.A(_05937_),
    .X(net241));
 sky130_fd_sc_hd__buf_4 fanout242 (.A(net248),
    .X(net242));
 sky130_fd_sc_hd__buf_4 fanout243 (.A(net248),
    .X(net243));
 sky130_fd_sc_hd__buf_4 fanout244 (.A(net248),
    .X(net244));
 sky130_fd_sc_hd__buf_4 fanout245 (.A(net248),
    .X(net245));
 sky130_fd_sc_hd__buf_4 fanout246 (.A(net248),
    .X(net246));
 sky130_fd_sc_hd__buf_8 fanout247 (.A(net248),
    .X(net247));
 sky130_fd_sc_hd__buf_6 fanout248 (.A(_05879_),
    .X(net248));
 sky130_fd_sc_hd__buf_4 fanout249 (.A(_05850_),
    .X(net249));
 sky130_fd_sc_hd__buf_4 fanout250 (.A(_05850_),
    .X(net250));
 sky130_fd_sc_hd__buf_2 fanout251 (.A(_05850_),
    .X(net251));
 sky130_fd_sc_hd__buf_6 fanout252 (.A(net253),
    .X(net252));
 sky130_fd_sc_hd__buf_6 fanout253 (.A(_05841_),
    .X(net253));
 sky130_fd_sc_hd__buf_6 fanout254 (.A(_05840_),
    .X(net254));
 sky130_fd_sc_hd__buf_12 fanout255 (.A(net257),
    .X(net255));
 sky130_fd_sc_hd__buf_8 fanout256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_16 fanout257 (.A(_02579_),
    .X(net257));
 sky130_fd_sc_hd__buf_4 fanout258 (.A(net259),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_8 fanout259 (.A(net261),
    .X(net259));
 sky130_fd_sc_hd__buf_8 fanout260 (.A(net261),
    .X(net260));
 sky130_fd_sc_hd__buf_12 fanout261 (.A(_02578_),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_4 fanout262 (.A(_08481_),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_2 fanout263 (.A(_08481_),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_4 fanout264 (.A(_08481_),
    .X(net264));
 sky130_fd_sc_hd__buf_2 fanout265 (.A(_08481_),
    .X(net265));
 sky130_fd_sc_hd__buf_8 fanout266 (.A(_06178_),
    .X(net266));
 sky130_fd_sc_hd__buf_2 fanout267 (.A(_06178_),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_4 fanout269 (.A(net270),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_4 fanout270 (.A(_05955_),
    .X(net270));
 sky130_fd_sc_hd__buf_4 fanout271 (.A(_05955_),
    .X(net271));
 sky130_fd_sc_hd__buf_4 fanout272 (.A(net276),
    .X(net272));
 sky130_fd_sc_hd__buf_6 fanout273 (.A(net275),
    .X(net273));
 sky130_fd_sc_hd__buf_6 fanout274 (.A(net275),
    .X(net274));
 sky130_fd_sc_hd__buf_4 fanout275 (.A(net276),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_4 fanout276 (.A(_05953_),
    .X(net276));
 sky130_fd_sc_hd__buf_6 fanout277 (.A(net279),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_4 fanout278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__buf_12 fanout279 (.A(_03357_),
    .X(net279));
 sky130_fd_sc_hd__buf_6 fanout280 (.A(net281),
    .X(net280));
 sky130_fd_sc_hd__buf_8 fanout281 (.A(_03346_),
    .X(net281));
 sky130_fd_sc_hd__buf_8 fanout282 (.A(_03291_),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_4 fanout283 (.A(net284),
    .X(net283));
 sky130_fd_sc_hd__buf_2 fanout284 (.A(net285),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_4 fanout285 (.A(net286),
    .X(net285));
 sky130_fd_sc_hd__buf_8 fanout286 (.A(_03247_),
    .X(net286));
 sky130_fd_sc_hd__buf_6 fanout287 (.A(net288),
    .X(net287));
 sky130_fd_sc_hd__buf_6 fanout288 (.A(net290),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_8 fanout289 (.A(net290),
    .X(net289));
 sky130_fd_sc_hd__buf_4 fanout290 (.A(net291),
    .X(net290));
 sky130_fd_sc_hd__buf_6 fanout291 (.A(net292),
    .X(net291));
 sky130_fd_sc_hd__buf_6 fanout292 (.A(_03236_),
    .X(net292));
 sky130_fd_sc_hd__buf_6 fanout293 (.A(net294),
    .X(net293));
 sky130_fd_sc_hd__buf_6 fanout294 (.A(net295),
    .X(net294));
 sky130_fd_sc_hd__buf_6 fanout295 (.A(net298),
    .X(net295));
 sky130_fd_sc_hd__buf_6 fanout296 (.A(net298),
    .X(net296));
 sky130_fd_sc_hd__buf_6 fanout297 (.A(net298),
    .X(net297));
 sky130_fd_sc_hd__buf_4 fanout298 (.A(_03225_),
    .X(net298));
 sky130_fd_sc_hd__buf_6 fanout299 (.A(_03225_),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_8 fanout300 (.A(net301),
    .X(net300));
 sky130_fd_sc_hd__buf_6 fanout301 (.A(net302),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_8 fanout302 (.A(net304),
    .X(net302));
 sky130_fd_sc_hd__buf_6 fanout303 (.A(net304),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_8 fanout304 (.A(_03214_),
    .X(net304));
 sky130_fd_sc_hd__buf_4 fanout305 (.A(net306),
    .X(net305));
 sky130_fd_sc_hd__buf_2 fanout306 (.A(net307),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_4 fanout307 (.A(net308),
    .X(net307));
 sky130_fd_sc_hd__buf_6 fanout308 (.A(net309),
    .X(net308));
 sky130_fd_sc_hd__buf_6 fanout309 (.A(_03203_),
    .X(net309));
 sky130_fd_sc_hd__buf_6 fanout310 (.A(\sel_op[2] ),
    .X(net310));
 sky130_fd_sc_hd__buf_6 fanout311 (.A(\sel_op[1] ),
    .X(net311));
 sky130_fd_sc_hd__buf_6 fanout312 (.A(net314),
    .X(net312));
 sky130_fd_sc_hd__buf_6 fanout313 (.A(net314),
    .X(net313));
 sky130_fd_sc_hd__buf_8 fanout314 (.A(\sel_op[0] ),
    .X(net314));
 sky130_fd_sc_hd__buf_8 fanout315 (.A(\op_code[3] ),
    .X(net315));
 sky130_fd_sc_hd__buf_6 fanout316 (.A(\op_code[2] ),
    .X(net316));
 sky130_fd_sc_hd__buf_6 fanout317 (.A(net325),
    .X(net317));
 sky130_fd_sc_hd__buf_8 fanout318 (.A(net324),
    .X(net318));
 sky130_fd_sc_hd__buf_8 fanout319 (.A(net324),
    .X(net319));
 sky130_fd_sc_hd__buf_2 fanout320 (.A(net324),
    .X(net320));
 sky130_fd_sc_hd__buf_6 fanout321 (.A(net324),
    .X(net321));
 sky130_fd_sc_hd__buf_2 fanout322 (.A(net324),
    .X(net322));
 sky130_fd_sc_hd__buf_6 fanout323 (.A(net324),
    .X(net323));
 sky130_fd_sc_hd__buf_12 fanout324 (.A(net325),
    .X(net324));
 sky130_fd_sc_hd__buf_8 fanout325 (.A(\cla_inst.in2[31] ),
    .X(net325));
 sky130_fd_sc_hd__buf_6 fanout326 (.A(net327),
    .X(net326));
 sky130_fd_sc_hd__buf_4 fanout327 (.A(\cla_inst.in2[30] ),
    .X(net327));
 sky130_fd_sc_hd__buf_6 fanout328 (.A(net334),
    .X(net328));
 sky130_fd_sc_hd__buf_6 fanout329 (.A(net330),
    .X(net329));
 sky130_fd_sc_hd__buf_6 fanout330 (.A(net334),
    .X(net330));
 sky130_fd_sc_hd__buf_6 fanout331 (.A(net332),
    .X(net331));
 sky130_fd_sc_hd__buf_4 fanout332 (.A(net334),
    .X(net332));
 sky130_fd_sc_hd__buf_6 fanout333 (.A(net334),
    .X(net333));
 sky130_fd_sc_hd__buf_6 fanout334 (.A(\cla_inst.in2[30] ),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_16 fanout335 (.A(\cla_inst.in2[29] ),
    .X(net335));
 sky130_fd_sc_hd__buf_6 fanout336 (.A(net337),
    .X(net336));
 sky130_fd_sc_hd__buf_8 fanout337 (.A(net339),
    .X(net337));
 sky130_fd_sc_hd__buf_12 fanout338 (.A(net339),
    .X(net338));
 sky130_fd_sc_hd__buf_8 fanout339 (.A(\cla_inst.in2[29] ),
    .X(net339));
 sky130_fd_sc_hd__buf_6 fanout340 (.A(net341),
    .X(net340));
 sky130_fd_sc_hd__buf_6 fanout341 (.A(net342),
    .X(net341));
 sky130_fd_sc_hd__buf_4 fanout342 (.A(\cla_inst.in2[28] ),
    .X(net342));
 sky130_fd_sc_hd__buf_6 fanout343 (.A(net344),
    .X(net343));
 sky130_fd_sc_hd__buf_8 fanout344 (.A(net348),
    .X(net344));
 sky130_fd_sc_hd__buf_8 fanout345 (.A(net346),
    .X(net345));
 sky130_fd_sc_hd__buf_12 fanout346 (.A(net348),
    .X(net346));
 sky130_fd_sc_hd__buf_4 fanout347 (.A(net348),
    .X(net347));
 sky130_fd_sc_hd__buf_8 fanout348 (.A(\cla_inst.in2[28] ),
    .X(net348));
 sky130_fd_sc_hd__buf_6 fanout349 (.A(net350),
    .X(net349));
 sky130_fd_sc_hd__buf_8 fanout350 (.A(net356),
    .X(net350));
 sky130_fd_sc_hd__buf_6 fanout351 (.A(net352),
    .X(net351));
 sky130_fd_sc_hd__buf_6 fanout352 (.A(net355),
    .X(net352));
 sky130_fd_sc_hd__buf_8 fanout353 (.A(net354),
    .X(net353));
 sky130_fd_sc_hd__buf_6 fanout354 (.A(net355),
    .X(net354));
 sky130_fd_sc_hd__buf_8 fanout355 (.A(net356),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_16 fanout356 (.A(\cla_inst.in2[27] ),
    .X(net356));
 sky130_fd_sc_hd__buf_8 fanout357 (.A(net358),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_16 fanout358 (.A(net362),
    .X(net358));
 sky130_fd_sc_hd__buf_12 fanout359 (.A(net362),
    .X(net359));
 sky130_fd_sc_hd__buf_6 fanout360 (.A(net361),
    .X(net360));
 sky130_fd_sc_hd__buf_6 fanout361 (.A(net362),
    .X(net361));
 sky130_fd_sc_hd__buf_12 fanout362 (.A(\cla_inst.in2[26] ),
    .X(net362));
 sky130_fd_sc_hd__buf_8 fanout363 (.A(net365),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_8 fanout364 (.A(net365),
    .X(net364));
 sky130_fd_sc_hd__buf_12 fanout365 (.A(net371),
    .X(net365));
 sky130_fd_sc_hd__buf_6 fanout366 (.A(net367),
    .X(net366));
 sky130_fd_sc_hd__buf_12 fanout367 (.A(net371),
    .X(net367));
 sky130_fd_sc_hd__buf_4 fanout368 (.A(net369),
    .X(net368));
 sky130_fd_sc_hd__buf_4 fanout369 (.A(net370),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_8 fanout370 (.A(net371),
    .X(net370));
 sky130_fd_sc_hd__buf_12 fanout371 (.A(\cla_inst.in2[25] ),
    .X(net371));
 sky130_fd_sc_hd__buf_8 fanout372 (.A(net374),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_8 fanout373 (.A(net374),
    .X(net373));
 sky130_fd_sc_hd__buf_12 fanout374 (.A(net380),
    .X(net374));
 sky130_fd_sc_hd__buf_6 fanout375 (.A(net376),
    .X(net375));
 sky130_fd_sc_hd__buf_12 fanout376 (.A(net380),
    .X(net376));
 sky130_fd_sc_hd__buf_6 fanout377 (.A(net379),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_8 fanout378 (.A(net379),
    .X(net378));
 sky130_fd_sc_hd__buf_4 fanout379 (.A(net380),
    .X(net379));
 sky130_fd_sc_hd__buf_12 fanout380 (.A(\cla_inst.in2[24] ),
    .X(net380));
 sky130_fd_sc_hd__buf_4 fanout381 (.A(net382),
    .X(net381));
 sky130_fd_sc_hd__buf_4 fanout382 (.A(\cla_inst.in2[23] ),
    .X(net382));
 sky130_fd_sc_hd__buf_6 fanout383 (.A(\cla_inst.in2[23] ),
    .X(net383));
 sky130_fd_sc_hd__buf_12 fanout384 (.A(net387),
    .X(net384));
 sky130_fd_sc_hd__buf_6 fanout385 (.A(net386),
    .X(net385));
 sky130_fd_sc_hd__buf_6 fanout386 (.A(net387),
    .X(net386));
 sky130_fd_sc_hd__buf_8 fanout387 (.A(\cla_inst.in2[23] ),
    .X(net387));
 sky130_fd_sc_hd__buf_6 fanout388 (.A(net389),
    .X(net388));
 sky130_fd_sc_hd__buf_8 fanout389 (.A(\cla_inst.in2[22] ),
    .X(net389));
 sky130_fd_sc_hd__buf_4 fanout390 (.A(net391),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_8 fanout391 (.A(\cla_inst.in2[22] ),
    .X(net391));
 sky130_fd_sc_hd__buf_8 fanout392 (.A(net393),
    .X(net392));
 sky130_fd_sc_hd__buf_8 fanout393 (.A(\cla_inst.in2[22] ),
    .X(net393));
 sky130_fd_sc_hd__buf_8 fanout394 (.A(net395),
    .X(net394));
 sky130_fd_sc_hd__buf_6 fanout395 (.A(\cla_inst.in2[22] ),
    .X(net395));
 sky130_fd_sc_hd__buf_8 fanout396 (.A(net399),
    .X(net396));
 sky130_fd_sc_hd__buf_6 fanout397 (.A(net398),
    .X(net397));
 sky130_fd_sc_hd__buf_6 fanout398 (.A(net399),
    .X(net398));
 sky130_fd_sc_hd__buf_8 fanout399 (.A(\cla_inst.in2[21] ),
    .X(net399));
 sky130_fd_sc_hd__buf_6 fanout400 (.A(net401),
    .X(net400));
 sky130_fd_sc_hd__buf_8 fanout401 (.A(net402),
    .X(net401));
 sky130_fd_sc_hd__buf_12 fanout402 (.A(\cla_inst.in2[21] ),
    .X(net402));
 sky130_fd_sc_hd__buf_4 fanout403 (.A(net404),
    .X(net403));
 sky130_fd_sc_hd__buf_6 fanout404 (.A(net405),
    .X(net404));
 sky130_fd_sc_hd__buf_4 fanout405 (.A(net406),
    .X(net405));
 sky130_fd_sc_hd__buf_8 fanout406 (.A(\cla_inst.in2[20] ),
    .X(net406));
 sky130_fd_sc_hd__buf_8 fanout407 (.A(\cla_inst.in2[20] ),
    .X(net407));
 sky130_fd_sc_hd__buf_6 fanout408 (.A(net409),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_4 fanout409 (.A(net410),
    .X(net409));
 sky130_fd_sc_hd__buf_8 fanout410 (.A(\cla_inst.in2[20] ),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_8 fanout411 (.A(net413),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_2 fanout412 (.A(net413),
    .X(net412));
 sky130_fd_sc_hd__buf_6 fanout413 (.A(net418),
    .X(net413));
 sky130_fd_sc_hd__buf_4 fanout414 (.A(net418),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_8 fanout415 (.A(net416),
    .X(net415));
 sky130_fd_sc_hd__buf_12 fanout416 (.A(net417),
    .X(net416));
 sky130_fd_sc_hd__buf_12 fanout417 (.A(net418),
    .X(net417));
 sky130_fd_sc_hd__buf_6 fanout418 (.A(\cla_inst.in2[19] ),
    .X(net418));
 sky130_fd_sc_hd__buf_6 fanout419 (.A(net420),
    .X(net419));
 sky130_fd_sc_hd__buf_6 fanout420 (.A(net421),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_8 fanout421 (.A(\cla_inst.in2[18] ),
    .X(net421));
 sky130_fd_sc_hd__buf_6 fanout422 (.A(\cla_inst.in2[18] ),
    .X(net422));
 sky130_fd_sc_hd__buf_6 fanout423 (.A(net425),
    .X(net423));
 sky130_fd_sc_hd__buf_6 fanout424 (.A(net425),
    .X(net424));
 sky130_fd_sc_hd__buf_8 fanout425 (.A(net426),
    .X(net425));
 sky130_fd_sc_hd__buf_6 fanout426 (.A(\cla_inst.in2[18] ),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_16 fanout427 (.A(net429),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_8 fanout428 (.A(net429),
    .X(net428));
 sky130_fd_sc_hd__buf_6 fanout429 (.A(net435),
    .X(net429));
 sky130_fd_sc_hd__buf_6 fanout430 (.A(net431),
    .X(net430));
 sky130_fd_sc_hd__buf_4 fanout431 (.A(net435),
    .X(net431));
 sky130_fd_sc_hd__buf_8 fanout432 (.A(net433),
    .X(net432));
 sky130_fd_sc_hd__buf_6 fanout433 (.A(net435),
    .X(net433));
 sky130_fd_sc_hd__buf_6 fanout434 (.A(net435),
    .X(net434));
 sky130_fd_sc_hd__buf_12 fanout435 (.A(\cla_inst.in2[17] ),
    .X(net435));
 sky130_fd_sc_hd__buf_6 fanout436 (.A(net437),
    .X(net436));
 sky130_fd_sc_hd__buf_8 fanout437 (.A(net438),
    .X(net437));
 sky130_fd_sc_hd__buf_6 fanout438 (.A(net441),
    .X(net438));
 sky130_fd_sc_hd__buf_8 fanout439 (.A(net441),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_4 fanout440 (.A(net441),
    .X(net440));
 sky130_fd_sc_hd__buf_8 fanout441 (.A(net445),
    .X(net441));
 sky130_fd_sc_hd__buf_6 fanout442 (.A(net443),
    .X(net442));
 sky130_fd_sc_hd__buf_4 fanout443 (.A(net444),
    .X(net443));
 sky130_fd_sc_hd__buf_12 fanout444 (.A(net445),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_16 fanout445 (.A(\cla_inst.in2[16] ),
    .X(net445));
 sky130_fd_sc_hd__buf_8 fanout446 (.A(net449),
    .X(net446));
 sky130_fd_sc_hd__buf_12 fanout447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__buf_12 fanout448 (.A(net449),
    .X(net448));
 sky130_fd_sc_hd__clkbuf_16 fanout449 (.A(\ApproximateM_inst.lob_16.lob2.genblk2.mux_final.sel ),
    .X(net449));
 sky130_fd_sc_hd__buf_12 fanout450 (.A(net453),
    .X(net450));
 sky130_fd_sc_hd__buf_6 fanout451 (.A(net452),
    .X(net451));
 sky130_fd_sc_hd__buf_8 fanout452 (.A(net453),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_16 fanout453 (.A(\ApproximateM_inst.lob_16.lob2.genblk2.mux_final.sel ),
    .X(net453));
 sky130_fd_sc_hd__buf_6 fanout454 (.A(net455),
    .X(net454));
 sky130_fd_sc_hd__buf_8 fanout455 (.A(net463),
    .X(net455));
 sky130_fd_sc_hd__buf_8 fanout456 (.A(net457),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_16 fanout457 (.A(net458),
    .X(net457));
 sky130_fd_sc_hd__buf_12 fanout458 (.A(net463),
    .X(net458));
 sky130_fd_sc_hd__buf_6 fanout459 (.A(net460),
    .X(net459));
 sky130_fd_sc_hd__buf_6 fanout460 (.A(net462),
    .X(net460));
 sky130_fd_sc_hd__buf_6 fanout461 (.A(net462),
    .X(net461));
 sky130_fd_sc_hd__buf_8 fanout462 (.A(net463),
    .X(net462));
 sky130_fd_sc_hd__clkbuf_16 fanout463 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[14].genblk1.mux.sel ),
    .X(net463));
 sky130_fd_sc_hd__buf_6 fanout464 (.A(net465),
    .X(net464));
 sky130_fd_sc_hd__buf_12 fanout465 (.A(net473),
    .X(net465));
 sky130_fd_sc_hd__buf_6 fanout466 (.A(net467),
    .X(net466));
 sky130_fd_sc_hd__clkbuf_16 fanout467 (.A(net468),
    .X(net467));
 sky130_fd_sc_hd__buf_6 fanout468 (.A(net473),
    .X(net468));
 sky130_fd_sc_hd__buf_6 fanout469 (.A(net470),
    .X(net469));
 sky130_fd_sc_hd__buf_4 fanout470 (.A(net472),
    .X(net470));
 sky130_fd_sc_hd__buf_6 fanout471 (.A(net472),
    .X(net471));
 sky130_fd_sc_hd__buf_8 fanout472 (.A(net473),
    .X(net472));
 sky130_fd_sc_hd__buf_8 fanout473 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[13].genblk1.mux.sel ),
    .X(net473));
 sky130_fd_sc_hd__buf_8 fanout474 (.A(net477),
    .X(net474));
 sky130_fd_sc_hd__buf_12 fanout475 (.A(net476),
    .X(net475));
 sky130_fd_sc_hd__buf_12 fanout476 (.A(net477),
    .X(net476));
 sky130_fd_sc_hd__buf_8 fanout477 (.A(net480),
    .X(net477));
 sky130_fd_sc_hd__buf_8 fanout478 (.A(net480),
    .X(net478));
 sky130_fd_sc_hd__buf_12 fanout479 (.A(net480),
    .X(net479));
 sky130_fd_sc_hd__clkbuf_16 fanout480 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[12].genblk1.mux.sel ),
    .X(net480));
 sky130_fd_sc_hd__clkbuf_8 fanout481 (.A(net482),
    .X(net481));
 sky130_fd_sc_hd__buf_4 fanout482 (.A(net483),
    .X(net482));
 sky130_fd_sc_hd__buf_6 fanout483 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[11].genblk1.mux.sel ),
    .X(net483));
 sky130_fd_sc_hd__buf_6 fanout484 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[11].genblk1.mux.sel ),
    .X(net484));
 sky130_fd_sc_hd__buf_2 fanout485 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[11].genblk1.mux.sel ),
    .X(net485));
 sky130_fd_sc_hd__buf_6 fanout486 (.A(net488),
    .X(net486));
 sky130_fd_sc_hd__buf_4 fanout487 (.A(net488),
    .X(net487));
 sky130_fd_sc_hd__buf_4 fanout488 (.A(net489),
    .X(net488));
 sky130_fd_sc_hd__buf_8 fanout489 (.A(net490),
    .X(net489));
 sky130_fd_sc_hd__buf_6 fanout490 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[11].genblk1.mux.sel ),
    .X(net490));
 sky130_fd_sc_hd__clkbuf_8 fanout491 (.A(net492),
    .X(net491));
 sky130_fd_sc_hd__buf_4 fanout492 (.A(net493),
    .X(net492));
 sky130_fd_sc_hd__buf_6 fanout493 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[10].genblk1.mux.sel ),
    .X(net493));
 sky130_fd_sc_hd__buf_6 fanout494 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[10].genblk1.mux.sel ),
    .X(net494));
 sky130_fd_sc_hd__buf_2 fanout495 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[10].genblk1.mux.sel ),
    .X(net495));
 sky130_fd_sc_hd__buf_8 fanout496 (.A(net498),
    .X(net496));
 sky130_fd_sc_hd__clkbuf_4 fanout497 (.A(net498),
    .X(net497));
 sky130_fd_sc_hd__buf_6 fanout498 (.A(net499),
    .X(net498));
 sky130_fd_sc_hd__buf_8 fanout499 (.A(net500),
    .X(net499));
 sky130_fd_sc_hd__buf_4 fanout500 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[10].genblk1.mux.sel ),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_4 fanout501 (.A(net502),
    .X(net501));
 sky130_fd_sc_hd__buf_6 fanout502 (.A(net503),
    .X(net502));
 sky130_fd_sc_hd__buf_8 fanout503 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[9].genblk1.mux.sel ),
    .X(net503));
 sky130_fd_sc_hd__buf_8 fanout504 (.A(net507),
    .X(net504));
 sky130_fd_sc_hd__buf_4 fanout505 (.A(net506),
    .X(net505));
 sky130_fd_sc_hd__buf_6 fanout506 (.A(net507),
    .X(net506));
 sky130_fd_sc_hd__clkbuf_16 fanout507 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[9].genblk1.mux.sel ),
    .X(net507));
 sky130_fd_sc_hd__clkbuf_8 fanout508 (.A(net509),
    .X(net508));
 sky130_fd_sc_hd__buf_4 fanout509 (.A(net510),
    .X(net509));
 sky130_fd_sc_hd__buf_6 fanout510 (.A(net511),
    .X(net510));
 sky130_fd_sc_hd__clkbuf_8 fanout511 (.A(net516),
    .X(net511));
 sky130_fd_sc_hd__buf_6 fanout512 (.A(net513),
    .X(net512));
 sky130_fd_sc_hd__buf_6 fanout513 (.A(net515),
    .X(net513));
 sky130_fd_sc_hd__buf_6 fanout514 (.A(net515),
    .X(net514));
 sky130_fd_sc_hd__buf_6 fanout515 (.A(net516),
    .X(net515));
 sky130_fd_sc_hd__buf_8 fanout516 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[8].genblk1.mux.sel ),
    .X(net516));
 sky130_fd_sc_hd__buf_6 fanout517 (.A(net518),
    .X(net517));
 sky130_fd_sc_hd__buf_6 fanout518 (.A(net519),
    .X(net518));
 sky130_fd_sc_hd__buf_8 fanout519 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[7].genblk1.mux.sel ),
    .X(net519));
 sky130_fd_sc_hd__buf_4 fanout520 (.A(net521),
    .X(net520));
 sky130_fd_sc_hd__buf_6 fanout521 (.A(net524),
    .X(net521));
 sky130_fd_sc_hd__buf_6 fanout522 (.A(net523),
    .X(net522));
 sky130_fd_sc_hd__buf_6 fanout523 (.A(net524),
    .X(net523));
 sky130_fd_sc_hd__buf_8 fanout524 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[7].genblk1.mux.sel ),
    .X(net524));
 sky130_fd_sc_hd__buf_4 fanout525 (.A(net527),
    .X(net525));
 sky130_fd_sc_hd__clkbuf_2 fanout526 (.A(net527),
    .X(net526));
 sky130_fd_sc_hd__buf_6 fanout527 (.A(net528),
    .X(net527));
 sky130_fd_sc_hd__clkbuf_4 fanout528 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[6].genblk1.mux.sel ),
    .X(net528));
 sky130_fd_sc_hd__clkbuf_8 fanout529 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[6].genblk1.mux.sel ),
    .X(net529));
 sky130_fd_sc_hd__buf_4 fanout530 (.A(net531),
    .X(net530));
 sky130_fd_sc_hd__buf_4 fanout531 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[6].genblk1.mux.sel ),
    .X(net531));
 sky130_fd_sc_hd__buf_8 fanout532 (.A(net534),
    .X(net532));
 sky130_fd_sc_hd__clkbuf_4 fanout533 (.A(net534),
    .X(net533));
 sky130_fd_sc_hd__buf_6 fanout534 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[6].genblk1.mux.sel ),
    .X(net534));
 sky130_fd_sc_hd__buf_6 fanout535 (.A(net536),
    .X(net535));
 sky130_fd_sc_hd__buf_6 fanout536 (.A(net549),
    .X(net536));
 sky130_fd_sc_hd__buf_6 fanout537 (.A(net539),
    .X(net537));
 sky130_fd_sc_hd__clkbuf_4 fanout538 (.A(net539),
    .X(net538));
 sky130_fd_sc_hd__buf_4 fanout539 (.A(net540),
    .X(net539));
 sky130_fd_sc_hd__buf_8 fanout540 (.A(net549),
    .X(net540));
 sky130_fd_sc_hd__buf_6 fanout541 (.A(net548),
    .X(net541));
 sky130_fd_sc_hd__buf_6 fanout542 (.A(net548),
    .X(net542));
 sky130_fd_sc_hd__buf_4 fanout543 (.A(net548),
    .X(net543));
 sky130_fd_sc_hd__clkbuf_8 fanout544 (.A(net548),
    .X(net544));
 sky130_fd_sc_hd__buf_4 fanout545 (.A(net547),
    .X(net545));
 sky130_fd_sc_hd__buf_4 fanout546 (.A(net547),
    .X(net546));
 sky130_fd_sc_hd__clkbuf_4 fanout547 (.A(net548),
    .X(net547));
 sky130_fd_sc_hd__buf_8 fanout548 (.A(net549),
    .X(net548));
 sky130_fd_sc_hd__buf_6 fanout549 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[5].genblk1.mux.sel ),
    .X(net549));
 sky130_fd_sc_hd__buf_6 fanout550 (.A(net551),
    .X(net550));
 sky130_fd_sc_hd__buf_6 fanout551 (.A(net563),
    .X(net551));
 sky130_fd_sc_hd__buf_6 fanout552 (.A(net554),
    .X(net552));
 sky130_fd_sc_hd__buf_4 fanout553 (.A(net554),
    .X(net553));
 sky130_fd_sc_hd__buf_6 fanout554 (.A(net563),
    .X(net554));
 sky130_fd_sc_hd__buf_6 fanout555 (.A(net563),
    .X(net555));
 sky130_fd_sc_hd__clkbuf_8 fanout556 (.A(net563),
    .X(net556));
 sky130_fd_sc_hd__buf_4 fanout557 (.A(net563),
    .X(net557));
 sky130_fd_sc_hd__buf_4 fanout558 (.A(net562),
    .X(net558));
 sky130_fd_sc_hd__buf_4 fanout559 (.A(net562),
    .X(net559));
 sky130_fd_sc_hd__buf_4 fanout560 (.A(net562),
    .X(net560));
 sky130_fd_sc_hd__buf_6 fanout561 (.A(net562),
    .X(net561));
 sky130_fd_sc_hd__buf_4 fanout562 (.A(net563),
    .X(net562));
 sky130_fd_sc_hd__buf_12 fanout563 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[4].genblk1.mux.sel ),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_8 fanout564 (.A(net565),
    .X(net564));
 sky130_fd_sc_hd__buf_8 fanout565 (.A(net571),
    .X(net565));
 sky130_fd_sc_hd__buf_6 fanout566 (.A(net567),
    .X(net566));
 sky130_fd_sc_hd__buf_8 fanout567 (.A(net571),
    .X(net567));
 sky130_fd_sc_hd__buf_4 fanout568 (.A(net571),
    .X(net568));
 sky130_fd_sc_hd__clkbuf_2 fanout569 (.A(net570),
    .X(net569));
 sky130_fd_sc_hd__buf_4 fanout570 (.A(net571),
    .X(net570));
 sky130_fd_sc_hd__clkbuf_8 fanout571 (.A(net580),
    .X(net571));
 sky130_fd_sc_hd__buf_4 fanout572 (.A(net580),
    .X(net572));
 sky130_fd_sc_hd__clkbuf_4 fanout573 (.A(net574),
    .X(net573));
 sky130_fd_sc_hd__buf_4 fanout574 (.A(net580),
    .X(net574));
 sky130_fd_sc_hd__clkbuf_8 fanout575 (.A(net576),
    .X(net575));
 sky130_fd_sc_hd__clkbuf_4 fanout576 (.A(net577),
    .X(net576));
 sky130_fd_sc_hd__buf_4 fanout577 (.A(net580),
    .X(net577));
 sky130_fd_sc_hd__buf_6 fanout578 (.A(net579),
    .X(net578));
 sky130_fd_sc_hd__buf_6 fanout579 (.A(net580),
    .X(net579));
 sky130_fd_sc_hd__buf_8 fanout580 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[3].genblk1.mux.sel ),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_4 fanout581 (.A(net582),
    .X(net581));
 sky130_fd_sc_hd__buf_2 fanout582 (.A(net586),
    .X(net582));
 sky130_fd_sc_hd__buf_6 fanout583 (.A(net586),
    .X(net583));
 sky130_fd_sc_hd__clkbuf_8 fanout584 (.A(net585),
    .X(net584));
 sky130_fd_sc_hd__buf_4 fanout585 (.A(net586),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_4 fanout586 (.A(net593),
    .X(net586));
 sky130_fd_sc_hd__buf_4 fanout587 (.A(net593),
    .X(net587));
 sky130_fd_sc_hd__buf_4 fanout588 (.A(net589),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_4 fanout589 (.A(net593),
    .X(net589));
 sky130_fd_sc_hd__clkbuf_8 fanout590 (.A(net591),
    .X(net590));
 sky130_fd_sc_hd__buf_6 fanout591 (.A(net592),
    .X(net591));
 sky130_fd_sc_hd__buf_4 fanout592 (.A(net593),
    .X(net592));
 sky130_fd_sc_hd__buf_4 fanout593 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[2].genblk1.mux.sel ),
    .X(net593));
 sky130_fd_sc_hd__buf_4 fanout594 (.A(net595),
    .X(net594));
 sky130_fd_sc_hd__buf_6 fanout595 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[1].genblk1.mux.sel ),
    .X(net595));
 sky130_fd_sc_hd__buf_4 fanout596 (.A(net597),
    .X(net596));
 sky130_fd_sc_hd__buf_6 fanout597 (.A(net598),
    .X(net597));
 sky130_fd_sc_hd__clkbuf_4 fanout598 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[1].genblk1.mux.sel ),
    .X(net598));
 sky130_fd_sc_hd__buf_2 fanout599 (.A(net600),
    .X(net599));
 sky130_fd_sc_hd__buf_4 fanout600 (.A(net605),
    .X(net600));
 sky130_fd_sc_hd__buf_4 fanout601 (.A(net605),
    .X(net601));
 sky130_fd_sc_hd__buf_4 fanout602 (.A(net604),
    .X(net602));
 sky130_fd_sc_hd__clkbuf_8 fanout603 (.A(net604),
    .X(net603));
 sky130_fd_sc_hd__buf_4 fanout604 (.A(net605),
    .X(net604));
 sky130_fd_sc_hd__clkbuf_8 fanout605 (.A(\ApproximateM_inst.lob_16.lob2.genblk1[1].genblk1.mux.sel ),
    .X(net605));
 sky130_fd_sc_hd__buf_4 fanout606 (.A(net608),
    .X(net606));
 sky130_fd_sc_hd__buf_4 fanout607 (.A(net608),
    .X(net607));
 sky130_fd_sc_hd__clkbuf_4 fanout608 (.A(net616),
    .X(net608));
 sky130_fd_sc_hd__buf_6 fanout609 (.A(net611),
    .X(net609));
 sky130_fd_sc_hd__clkbuf_4 fanout610 (.A(net611),
    .X(net610));
 sky130_fd_sc_hd__clkbuf_8 fanout611 (.A(net616),
    .X(net611));
 sky130_fd_sc_hd__buf_4 fanout612 (.A(net614),
    .X(net612));
 sky130_fd_sc_hd__clkbuf_4 fanout613 (.A(net614),
    .X(net613));
 sky130_fd_sc_hd__buf_6 fanout614 (.A(net616),
    .X(net614));
 sky130_fd_sc_hd__buf_6 fanout615 (.A(net616),
    .X(net615));
 sky130_fd_sc_hd__buf_4 fanout616 (.A(\ApproximateM_inst.lob_16.lob2.mux.sel ),
    .X(net616));
 sky130_fd_sc_hd__buf_6 fanout617 (.A(net618),
    .X(net617));
 sky130_fd_sc_hd__buf_8 fanout618 (.A(\cla_inst.in1[31] ),
    .X(net618));
 sky130_fd_sc_hd__buf_6 fanout619 (.A(net624),
    .X(net619));
 sky130_fd_sc_hd__buf_4 fanout620 (.A(net621),
    .X(net620));
 sky130_fd_sc_hd__buf_4 fanout621 (.A(net624),
    .X(net621));
 sky130_fd_sc_hd__buf_6 fanout622 (.A(net624),
    .X(net622));
 sky130_fd_sc_hd__buf_4 fanout623 (.A(net624),
    .X(net623));
 sky130_fd_sc_hd__buf_6 fanout624 (.A(\cla_inst.in1[31] ),
    .X(net624));
 sky130_fd_sc_hd__buf_8 fanout625 (.A(net626),
    .X(net625));
 sky130_fd_sc_hd__buf_6 fanout626 (.A(\cla_inst.in1[30] ),
    .X(net626));
 sky130_fd_sc_hd__buf_6 fanout627 (.A(net632),
    .X(net627));
 sky130_fd_sc_hd__buf_6 fanout628 (.A(net629),
    .X(net628));
 sky130_fd_sc_hd__clkbuf_4 fanout629 (.A(net632),
    .X(net629));
 sky130_fd_sc_hd__buf_6 fanout630 (.A(net631),
    .X(net630));
 sky130_fd_sc_hd__buf_6 fanout631 (.A(net632),
    .X(net631));
 sky130_fd_sc_hd__buf_6 fanout632 (.A(\cla_inst.in1[30] ),
    .X(net632));
 sky130_fd_sc_hd__buf_8 fanout633 (.A(net634),
    .X(net633));
 sky130_fd_sc_hd__buf_8 fanout634 (.A(\cla_inst.in1[29] ),
    .X(net634));
 sky130_fd_sc_hd__buf_6 fanout635 (.A(net641),
    .X(net635));
 sky130_fd_sc_hd__clkbuf_4 fanout636 (.A(net641),
    .X(net636));
 sky130_fd_sc_hd__buf_4 fanout637 (.A(net641),
    .X(net637));
 sky130_fd_sc_hd__buf_2 fanout638 (.A(net641),
    .X(net638));
 sky130_fd_sc_hd__buf_6 fanout639 (.A(net640),
    .X(net639));
 sky130_fd_sc_hd__buf_8 fanout640 (.A(net641),
    .X(net640));
 sky130_fd_sc_hd__buf_6 fanout641 (.A(\cla_inst.in1[29] ),
    .X(net641));
 sky130_fd_sc_hd__buf_8 fanout642 (.A(net643),
    .X(net642));
 sky130_fd_sc_hd__buf_6 fanout643 (.A(\cla_inst.in1[28] ),
    .X(net643));
 sky130_fd_sc_hd__buf_6 fanout644 (.A(net645),
    .X(net644));
 sky130_fd_sc_hd__buf_8 fanout645 (.A(\cla_inst.in1[28] ),
    .X(net645));
 sky130_fd_sc_hd__clkbuf_8 fanout646 (.A(net650),
    .X(net646));
 sky130_fd_sc_hd__buf_2 fanout647 (.A(net650),
    .X(net647));
 sky130_fd_sc_hd__buf_6 fanout648 (.A(net649),
    .X(net648));
 sky130_fd_sc_hd__buf_6 fanout649 (.A(net650),
    .X(net649));
 sky130_fd_sc_hd__buf_6 fanout650 (.A(\cla_inst.in1[28] ),
    .X(net650));
 sky130_fd_sc_hd__buf_6 fanout651 (.A(net652),
    .X(net651));
 sky130_fd_sc_hd__buf_4 fanout652 (.A(net653),
    .X(net652));
 sky130_fd_sc_hd__buf_4 fanout653 (.A(\cla_inst.in1[27] ),
    .X(net653));
 sky130_fd_sc_hd__buf_6 fanout654 (.A(net655),
    .X(net654));
 sky130_fd_sc_hd__clkbuf_16 fanout655 (.A(\cla_inst.in1[27] ),
    .X(net655));
 sky130_fd_sc_hd__buf_6 fanout656 (.A(net657),
    .X(net656));
 sky130_fd_sc_hd__buf_8 fanout657 (.A(net658),
    .X(net657));
 sky130_fd_sc_hd__buf_6 fanout658 (.A(\cla_inst.in1[27] ),
    .X(net658));
 sky130_fd_sc_hd__buf_4 fanout659 (.A(net660),
    .X(net659));
 sky130_fd_sc_hd__buf_4 fanout660 (.A(net661),
    .X(net660));
 sky130_fd_sc_hd__buf_6 fanout661 (.A(\cla_inst.in1[26] ),
    .X(net661));
 sky130_fd_sc_hd__buf_6 fanout662 (.A(net663),
    .X(net662));
 sky130_fd_sc_hd__buf_12 fanout663 (.A(\cla_inst.in1[26] ),
    .X(net663));
 sky130_fd_sc_hd__buf_6 fanout664 (.A(net665),
    .X(net664));
 sky130_fd_sc_hd__buf_6 fanout665 (.A(net666),
    .X(net665));
 sky130_fd_sc_hd__buf_4 fanout666 (.A(\cla_inst.in1[26] ),
    .X(net666));
 sky130_fd_sc_hd__buf_4 fanout667 (.A(net668),
    .X(net667));
 sky130_fd_sc_hd__buf_8 fanout668 (.A(net669),
    .X(net668));
 sky130_fd_sc_hd__buf_6 fanout669 (.A(net675),
    .X(net669));
 sky130_fd_sc_hd__buf_8 fanout670 (.A(net671),
    .X(net670));
 sky130_fd_sc_hd__buf_6 fanout671 (.A(net675),
    .X(net671));
 sky130_fd_sc_hd__buf_6 fanout672 (.A(net674),
    .X(net672));
 sky130_fd_sc_hd__clkbuf_4 fanout673 (.A(net674),
    .X(net673));
 sky130_fd_sc_hd__buf_8 fanout674 (.A(net675),
    .X(net674));
 sky130_fd_sc_hd__buf_6 fanout675 (.A(\cla_inst.in1[25] ),
    .X(net675));
 sky130_fd_sc_hd__buf_6 fanout676 (.A(net677),
    .X(net676));
 sky130_fd_sc_hd__buf_8 fanout677 (.A(net679),
    .X(net677));
 sky130_fd_sc_hd__buf_6 fanout678 (.A(net679),
    .X(net678));
 sky130_fd_sc_hd__buf_6 fanout679 (.A(\cla_inst.in1[24] ),
    .X(net679));
 sky130_fd_sc_hd__buf_8 fanout680 (.A(net683),
    .X(net680));
 sky130_fd_sc_hd__buf_8 fanout681 (.A(net683),
    .X(net681));
 sky130_fd_sc_hd__buf_4 fanout682 (.A(net683),
    .X(net682));
 sky130_fd_sc_hd__buf_6 fanout683 (.A(net684),
    .X(net683));
 sky130_fd_sc_hd__buf_4 fanout684 (.A(\cla_inst.in1[24] ),
    .X(net684));
 sky130_fd_sc_hd__clkbuf_8 fanout685 (.A(net686),
    .X(net685));
 sky130_fd_sc_hd__buf_12 fanout686 (.A(net693),
    .X(net686));
 sky130_fd_sc_hd__buf_6 fanout687 (.A(net688),
    .X(net687));
 sky130_fd_sc_hd__clkbuf_8 fanout688 (.A(net693),
    .X(net688));
 sky130_fd_sc_hd__clkbuf_16 fanout689 (.A(net693),
    .X(net689));
 sky130_fd_sc_hd__buf_8 fanout690 (.A(net693),
    .X(net690));
 sky130_fd_sc_hd__buf_6 fanout691 (.A(net692),
    .X(net691));
 sky130_fd_sc_hd__buf_4 fanout692 (.A(net693),
    .X(net692));
 sky130_fd_sc_hd__buf_8 fanout693 (.A(\cla_inst.in1[23] ),
    .X(net693));
 sky130_fd_sc_hd__buf_6 fanout694 (.A(net695),
    .X(net694));
 sky130_fd_sc_hd__buf_8 fanout695 (.A(net701),
    .X(net695));
 sky130_fd_sc_hd__buf_4 fanout696 (.A(net697),
    .X(net696));
 sky130_fd_sc_hd__buf_4 fanout697 (.A(net701),
    .X(net697));
 sky130_fd_sc_hd__clkbuf_16 fanout698 (.A(net699),
    .X(net698));
 sky130_fd_sc_hd__clkbuf_16 fanout699 (.A(net700),
    .X(net699));
 sky130_fd_sc_hd__buf_12 fanout700 (.A(net701),
    .X(net700));
 sky130_fd_sc_hd__clkbuf_16 fanout701 (.A(\cla_inst.in1[22] ),
    .X(net701));
 sky130_fd_sc_hd__buf_6 fanout702 (.A(net703),
    .X(net702));
 sky130_fd_sc_hd__buf_8 fanout703 (.A(net710),
    .X(net703));
 sky130_fd_sc_hd__buf_6 fanout704 (.A(net710),
    .X(net704));
 sky130_fd_sc_hd__buf_2 fanout705 (.A(net710),
    .X(net705));
 sky130_fd_sc_hd__buf_8 fanout706 (.A(net708),
    .X(net706));
 sky130_fd_sc_hd__buf_8 fanout707 (.A(net708),
    .X(net707));
 sky130_fd_sc_hd__buf_8 fanout708 (.A(net710),
    .X(net708));
 sky130_fd_sc_hd__buf_6 fanout709 (.A(net710),
    .X(net709));
 sky130_fd_sc_hd__buf_12 fanout710 (.A(\cla_inst.in1[21] ),
    .X(net710));
 sky130_fd_sc_hd__clkbuf_8 fanout711 (.A(net712),
    .X(net711));
 sky130_fd_sc_hd__buf_6 fanout712 (.A(net719),
    .X(net712));
 sky130_fd_sc_hd__buf_6 fanout713 (.A(net714),
    .X(net713));
 sky130_fd_sc_hd__clkbuf_8 fanout714 (.A(net719),
    .X(net714));
 sky130_fd_sc_hd__buf_8 fanout715 (.A(net718),
    .X(net715));
 sky130_fd_sc_hd__buf_4 fanout716 (.A(net718),
    .X(net716));
 sky130_fd_sc_hd__buf_6 fanout717 (.A(net718),
    .X(net717));
 sky130_fd_sc_hd__buf_8 fanout718 (.A(net719),
    .X(net718));
 sky130_fd_sc_hd__buf_6 fanout719 (.A(\cla_inst.in1[20] ),
    .X(net719));
 sky130_fd_sc_hd__buf_6 fanout720 (.A(net721),
    .X(net720));
 sky130_fd_sc_hd__buf_8 fanout721 (.A(net724),
    .X(net721));
 sky130_fd_sc_hd__buf_4 fanout722 (.A(net723),
    .X(net722));
 sky130_fd_sc_hd__clkbuf_8 fanout723 (.A(net724),
    .X(net723));
 sky130_fd_sc_hd__buf_6 fanout724 (.A(\cla_inst.in1[19] ),
    .X(net724));
 sky130_fd_sc_hd__buf_6 fanout725 (.A(net728),
    .X(net725));
 sky130_fd_sc_hd__buf_6 fanout726 (.A(net728),
    .X(net726));
 sky130_fd_sc_hd__buf_8 fanout727 (.A(net728),
    .X(net727));
 sky130_fd_sc_hd__buf_12 fanout728 (.A(\cla_inst.in1[19] ),
    .X(net728));
 sky130_fd_sc_hd__buf_6 fanout729 (.A(net730),
    .X(net729));
 sky130_fd_sc_hd__buf_12 fanout730 (.A(net736),
    .X(net730));
 sky130_fd_sc_hd__buf_4 fanout731 (.A(net732),
    .X(net731));
 sky130_fd_sc_hd__buf_6 fanout732 (.A(net736),
    .X(net732));
 sky130_fd_sc_hd__buf_8 fanout733 (.A(net735),
    .X(net733));
 sky130_fd_sc_hd__buf_8 fanout734 (.A(net735),
    .X(net734));
 sky130_fd_sc_hd__buf_12 fanout735 (.A(net736),
    .X(net735));
 sky130_fd_sc_hd__buf_12 fanout736 (.A(\cla_inst.in1[18] ),
    .X(net736));
 sky130_fd_sc_hd__buf_6 fanout737 (.A(net739),
    .X(net737));
 sky130_fd_sc_hd__buf_8 fanout738 (.A(net739),
    .X(net738));
 sky130_fd_sc_hd__clkbuf_8 fanout739 (.A(net745),
    .X(net739));
 sky130_fd_sc_hd__buf_4 fanout740 (.A(net741),
    .X(net740));
 sky130_fd_sc_hd__buf_6 fanout741 (.A(net745),
    .X(net741));
 sky130_fd_sc_hd__buf_12 fanout742 (.A(net744),
    .X(net742));
 sky130_fd_sc_hd__buf_8 fanout743 (.A(net744),
    .X(net743));
 sky130_fd_sc_hd__clkbuf_16 fanout744 (.A(net745),
    .X(net744));
 sky130_fd_sc_hd__buf_8 fanout745 (.A(\cla_inst.in1[17] ),
    .X(net745));
 sky130_fd_sc_hd__buf_12 fanout746 (.A(net754),
    .X(net746));
 sky130_fd_sc_hd__buf_8 fanout747 (.A(net754),
    .X(net747));
 sky130_fd_sc_hd__buf_4 fanout748 (.A(net749),
    .X(net748));
 sky130_fd_sc_hd__buf_6 fanout749 (.A(net750),
    .X(net749));
 sky130_fd_sc_hd__buf_4 fanout750 (.A(net754),
    .X(net750));
 sky130_fd_sc_hd__buf_12 fanout751 (.A(net753),
    .X(net751));
 sky130_fd_sc_hd__clkbuf_8 fanout752 (.A(net753),
    .X(net752));
 sky130_fd_sc_hd__clkbuf_16 fanout753 (.A(net754),
    .X(net753));
 sky130_fd_sc_hd__buf_8 fanout754 (.A(\cla_inst.in1[16] ),
    .X(net754));
 sky130_fd_sc_hd__buf_8 fanout755 (.A(net756),
    .X(net755));
 sky130_fd_sc_hd__buf_8 fanout756 (.A(net760),
    .X(net756));
 sky130_fd_sc_hd__buf_4 fanout757 (.A(net759),
    .X(net757));
 sky130_fd_sc_hd__clkbuf_4 fanout758 (.A(net759),
    .X(net758));
 sky130_fd_sc_hd__buf_8 fanout759 (.A(net760),
    .X(net759));
 sky130_fd_sc_hd__buf_6 fanout760 (.A(\ApproximateM_inst.lob_16.lob1.genblk2.mux_final.sel ),
    .X(net760));
 sky130_fd_sc_hd__buf_8 fanout761 (.A(net765),
    .X(net761));
 sky130_fd_sc_hd__buf_4 fanout762 (.A(net763),
    .X(net762));
 sky130_fd_sc_hd__buf_6 fanout763 (.A(net764),
    .X(net763));
 sky130_fd_sc_hd__buf_6 fanout764 (.A(net765),
    .X(net764));
 sky130_fd_sc_hd__buf_12 fanout765 (.A(\ApproximateM_inst.lob_16.lob1.genblk2.mux_final.sel ),
    .X(net765));
 sky130_fd_sc_hd__buf_12 fanout766 (.A(net772),
    .X(net766));
 sky130_fd_sc_hd__buf_6 fanout767 (.A(net772),
    .X(net767));
 sky130_fd_sc_hd__buf_4 fanout768 (.A(net769),
    .X(net768));
 sky130_fd_sc_hd__clkbuf_4 fanout769 (.A(net770),
    .X(net769));
 sky130_fd_sc_hd__buf_6 fanout770 (.A(net772),
    .X(net770));
 sky130_fd_sc_hd__buf_12 fanout771 (.A(net772),
    .X(net771));
 sky130_fd_sc_hd__buf_12 fanout772 (.A(\ApproximateM_inst.lob_16.lob1.genblk1[14].genblk1.mux.sel ),
    .X(net772));
 sky130_fd_sc_hd__buf_6 fanout773 (.A(net776),
    .X(net773));
 sky130_fd_sc_hd__buf_6 fanout774 (.A(net775),
    .X(net774));
 sky130_fd_sc_hd__buf_4 fanout775 (.A(net776),
    .X(net775));
 sky130_fd_sc_hd__buf_12 fanout776 (.A(\ApproximateM_inst.lob_16.lob1.genblk1[14].genblk1.mux.sel ),
    .X(net776));
 sky130_fd_sc_hd__buf_6 fanout777 (.A(net778),
    .X(net777));
 sky130_fd_sc_hd__clkbuf_16 fanout778 (.A(net787),
    .X(net778));
 sky130_fd_sc_hd__buf_8 fanout779 (.A(net787),
    .X(net779));
 sky130_fd_sc_hd__clkbuf_16 fanout780 (.A(net783),
    .X(net780));
 sky130_fd_sc_hd__buf_6 fanout781 (.A(net782),
    .X(net781));
 sky130_fd_sc_hd__buf_8 fanout782 (.A(net783),
    .X(net782));
 sky130_fd_sc_hd__buf_4 fanout783 (.A(net787),
    .X(net783));
 sky130_fd_sc_hd__buf_6 fanout784 (.A(net785),
    .X(net784));
 sky130_fd_sc_hd__clkbuf_8 fanout785 (.A(net786),
    .X(net785));
 sky130_fd_sc_hd__clkbuf_2 fanout786 (.A(net787),
    .X(net786));
 sky130_fd_sc_hd__buf_12 fanout787 (.A(\ApproximateM_inst.lob_16.lob1.genblk1[13].genblk1.mux.sel ),
    .X(net787));
 sky130_fd_sc_hd__buf_6 fanout788 (.A(net789),
    .X(net788));
 sky130_fd_sc_hd__buf_6 fanout789 (.A(net790),
    .X(net789));
 sky130_fd_sc_hd__buf_6 fanout790 (.A(net799),
    .X(net790));
 sky130_fd_sc_hd__clkbuf_8 fanout791 (.A(net794),
    .X(net791));
 sky130_fd_sc_hd__buf_6 fanout792 (.A(net793),
    .X(net792));
 sky130_fd_sc_hd__buf_12 fanout793 (.A(net794),
    .X(net793));
 sky130_fd_sc_hd__buf_6 fanout794 (.A(net799),
    .X(net794));
 sky130_fd_sc_hd__buf_8 fanout795 (.A(net799),
    .X(net795));
 sky130_fd_sc_hd__clkbuf_8 fanout796 (.A(net798),
    .X(net796));
 sky130_fd_sc_hd__buf_12 fanout797 (.A(net798),
    .X(net797));
 sky130_fd_sc_hd__buf_6 fanout798 (.A(net799),
    .X(net798));
 sky130_fd_sc_hd__buf_8 fanout799 (.A(\ApproximateM_inst.lob_16.lob1.genblk1[12].genblk1.mux.sel ),
    .X(net799));
 sky130_fd_sc_hd__clkbuf_16 fanout800 (.A(net803),
    .X(net800));
 sky130_fd_sc_hd__buf_6 fanout801 (.A(net803),
    .X(net801));
 sky130_fd_sc_hd__buf_8 fanout802 (.A(net803),
    .X(net802));
 sky130_fd_sc_hd__buf_6 fanout803 (.A(net809),
    .X(net803));
 sky130_fd_sc_hd__buf_4 fanout804 (.A(net809),
    .X(net804));
 sky130_fd_sc_hd__buf_6 fanout805 (.A(net806),
    .X(net805));
 sky130_fd_sc_hd__clkbuf_16 fanout806 (.A(net809),
    .X(net806));
 sky130_fd_sc_hd__buf_6 fanout807 (.A(net809),
    .X(net807));
 sky130_fd_sc_hd__buf_6 fanout808 (.A(net809),
    .X(net808));
 sky130_fd_sc_hd__buf_8 fanout809 (.A(\ApproximateM_inst.lob_16.lob1.genblk1[11].genblk1.mux.sel ),
    .X(net809));
 sky130_fd_sc_hd__buf_12 fanout810 (.A(net813),
    .X(net810));
 sky130_fd_sc_hd__buf_4 fanout811 (.A(net813),
    .X(net811));
 sky130_fd_sc_hd__buf_6 fanout812 (.A(net813),
    .X(net812));
 sky130_fd_sc_hd__buf_6 fanout813 (.A(\ApproximateM_inst.lob_16.lob1.genblk1[10].genblk1.mux.sel ),
    .X(net813));
 sky130_fd_sc_hd__buf_6 fanout814 (.A(net815),
    .X(net814));
 sky130_fd_sc_hd__buf_12 fanout815 (.A(net820),
    .X(net815));
 sky130_fd_sc_hd__clkbuf_8 fanout816 (.A(net818),
    .X(net816));
 sky130_fd_sc_hd__clkbuf_2 fanout817 (.A(net818),
    .X(net817));
 sky130_fd_sc_hd__buf_6 fanout818 (.A(net819),
    .X(net818));
 sky130_fd_sc_hd__clkbuf_4 fanout819 (.A(net820),
    .X(net819));
 sky130_fd_sc_hd__buf_6 fanout820 (.A(\ApproximateM_inst.lob_16.lob1.genblk1[10].genblk1.mux.sel ),
    .X(net820));
 sky130_fd_sc_hd__buf_8 fanout821 (.A(net824),
    .X(net821));
 sky130_fd_sc_hd__buf_4 fanout822 (.A(net824),
    .X(net822));
 sky130_fd_sc_hd__clkbuf_16 fanout823 (.A(net824),
    .X(net823));
 sky130_fd_sc_hd__buf_6 fanout824 (.A(\ApproximateM_inst.lob_16.lob1.genblk1[9].genblk1.mux.sel ),
    .X(net824));
 sky130_fd_sc_hd__buf_6 fanout825 (.A(net826),
    .X(net825));
 sky130_fd_sc_hd__buf_8 fanout826 (.A(\ApproximateM_inst.lob_16.lob1.genblk1[9].genblk1.mux.sel ),
    .X(net826));
 sky130_fd_sc_hd__buf_8 fanout827 (.A(net828),
    .X(net827));
 sky130_fd_sc_hd__buf_6 fanout828 (.A(net829),
    .X(net828));
 sky130_fd_sc_hd__buf_6 fanout829 (.A(\ApproximateM_inst.lob_16.lob1.genblk1[9].genblk1.mux.sel ),
    .X(net829));
 sky130_fd_sc_hd__buf_6 fanout830 (.A(net832),
    .X(net830));
 sky130_fd_sc_hd__buf_8 fanout831 (.A(net832),
    .X(net831));
 sky130_fd_sc_hd__buf_12 fanout832 (.A(net839),
    .X(net832));
 sky130_fd_sc_hd__buf_12 fanout833 (.A(net839),
    .X(net833));
 sky130_fd_sc_hd__clkbuf_4 fanout834 (.A(net839),
    .X(net834));
 sky130_fd_sc_hd__clkbuf_8 fanout835 (.A(net836),
    .X(net835));
 sky130_fd_sc_hd__clkbuf_8 fanout836 (.A(net837),
    .X(net836));
 sky130_fd_sc_hd__buf_6 fanout837 (.A(net839),
    .X(net837));
 sky130_fd_sc_hd__clkbuf_8 fanout838 (.A(net839),
    .X(net838));
 sky130_fd_sc_hd__buf_12 fanout839 (.A(\ApproximateM_inst.lob_16.lob1.genblk1[8].genblk1.mux.sel ),
    .X(net839));
 sky130_fd_sc_hd__buf_8 fanout840 (.A(net842),
    .X(net840));
 sky130_fd_sc_hd__buf_8 fanout841 (.A(net842),
    .X(net841));
 sky130_fd_sc_hd__buf_12 fanout842 (.A(\ApproximateM_inst.lob_16.lob1.genblk1[7].genblk1.mux.sel ),
    .X(net842));
 sky130_fd_sc_hd__buf_12 fanout843 (.A(net849),
    .X(net843));
 sky130_fd_sc_hd__buf_6 fanout844 (.A(net849),
    .X(net844));
 sky130_fd_sc_hd__buf_6 fanout845 (.A(net849),
    .X(net845));
 sky130_fd_sc_hd__buf_6 fanout846 (.A(net847),
    .X(net846));
 sky130_fd_sc_hd__buf_4 fanout847 (.A(net848),
    .X(net847));
 sky130_fd_sc_hd__buf_6 fanout848 (.A(net849),
    .X(net848));
 sky130_fd_sc_hd__buf_8 fanout849 (.A(\ApproximateM_inst.lob_16.lob1.genblk1[7].genblk1.mux.sel ),
    .X(net849));
 sky130_fd_sc_hd__buf_6 fanout850 (.A(net852),
    .X(net850));
 sky130_fd_sc_hd__buf_2 fanout851 (.A(net852),
    .X(net851));
 sky130_fd_sc_hd__buf_12 fanout852 (.A(\ApproximateM_inst.lob_16.lob1.genblk1[6].genblk1.mux.sel ),
    .X(net852));
 sky130_fd_sc_hd__clkbuf_16 fanout853 (.A(net854),
    .X(net853));
 sky130_fd_sc_hd__buf_12 fanout854 (.A(net859),
    .X(net854));
 sky130_fd_sc_hd__clkbuf_8 fanout855 (.A(net859),
    .X(net855));
 sky130_fd_sc_hd__buf_8 fanout856 (.A(net857),
    .X(net856));
 sky130_fd_sc_hd__buf_6 fanout857 (.A(net858),
    .X(net857));
 sky130_fd_sc_hd__buf_6 fanout858 (.A(net859),
    .X(net858));
 sky130_fd_sc_hd__buf_12 fanout859 (.A(\ApproximateM_inst.lob_16.lob1.genblk1[6].genblk1.mux.sel ),
    .X(net859));
 sky130_fd_sc_hd__buf_6 fanout860 (.A(net862),
    .X(net860));
 sky130_fd_sc_hd__buf_6 fanout861 (.A(net862),
    .X(net861));
 sky130_fd_sc_hd__buf_6 fanout862 (.A(net869),
    .X(net862));
 sky130_fd_sc_hd__buf_8 fanout863 (.A(net864),
    .X(net863));
 sky130_fd_sc_hd__buf_12 fanout864 (.A(net869),
    .X(net864));
 sky130_fd_sc_hd__clkbuf_8 fanout865 (.A(net867),
    .X(net865));
 sky130_fd_sc_hd__buf_6 fanout866 (.A(net867),
    .X(net866));
 sky130_fd_sc_hd__buf_6 fanout867 (.A(net868),
    .X(net867));
 sky130_fd_sc_hd__clkbuf_8 fanout868 (.A(net869),
    .X(net868));
 sky130_fd_sc_hd__buf_12 fanout869 (.A(\ApproximateM_inst.lob_16.lob1.genblk1[5].genblk1.mux.sel ),
    .X(net869));
 sky130_fd_sc_hd__buf_6 fanout870 (.A(net871),
    .X(net870));
 sky130_fd_sc_hd__buf_8 fanout871 (.A(net879),
    .X(net871));
 sky130_fd_sc_hd__buf_6 fanout872 (.A(net874),
    .X(net872));
 sky130_fd_sc_hd__buf_8 fanout873 (.A(net874),
    .X(net873));
 sky130_fd_sc_hd__buf_12 fanout874 (.A(net879),
    .X(net874));
 sky130_fd_sc_hd__clkbuf_8 fanout875 (.A(net878),
    .X(net875));
 sky130_fd_sc_hd__buf_6 fanout876 (.A(net877),
    .X(net876));
 sky130_fd_sc_hd__buf_6 fanout877 (.A(net878),
    .X(net877));
 sky130_fd_sc_hd__clkbuf_8 fanout878 (.A(net879),
    .X(net878));
 sky130_fd_sc_hd__clkbuf_16 fanout879 (.A(\ApproximateM_inst.lob_16.lob1.genblk1[4].genblk1.mux.sel ),
    .X(net879));
 sky130_fd_sc_hd__buf_6 fanout880 (.A(net891),
    .X(net880));
 sky130_fd_sc_hd__clkbuf_4 fanout881 (.A(net891),
    .X(net881));
 sky130_fd_sc_hd__buf_4 fanout882 (.A(net885),
    .X(net882));
 sky130_fd_sc_hd__buf_8 fanout883 (.A(net885),
    .X(net883));
 sky130_fd_sc_hd__clkbuf_4 fanout884 (.A(net885),
    .X(net884));
 sky130_fd_sc_hd__buf_6 fanout885 (.A(net891),
    .X(net885));
 sky130_fd_sc_hd__clkbuf_8 fanout886 (.A(net890),
    .X(net886));
 sky130_fd_sc_hd__buf_6 fanout887 (.A(net889),
    .X(net887));
 sky130_fd_sc_hd__buf_2 fanout888 (.A(net889),
    .X(net888));
 sky130_fd_sc_hd__buf_8 fanout889 (.A(net890),
    .X(net889));
 sky130_fd_sc_hd__buf_4 fanout890 (.A(net891),
    .X(net890));
 sky130_fd_sc_hd__buf_12 fanout891 (.A(\ApproximateM_inst.lob_16.lob1.genblk1[3].genblk1.mux.sel ),
    .X(net891));
 sky130_fd_sc_hd__buf_4 fanout892 (.A(net893),
    .X(net892));
 sky130_fd_sc_hd__buf_8 fanout893 (.A(net896),
    .X(net893));
 sky130_fd_sc_hd__buf_6 fanout894 (.A(net895),
    .X(net894));
 sky130_fd_sc_hd__buf_8 fanout895 (.A(net896),
    .X(net895));
 sky130_fd_sc_hd__buf_8 fanout896 (.A(\ApproximateM_inst.lob_16.lob1.genblk1[2].genblk1.mux.sel ),
    .X(net896));
 sky130_fd_sc_hd__clkbuf_8 fanout897 (.A(net898),
    .X(net897));
 sky130_fd_sc_hd__buf_4 fanout898 (.A(net900),
    .X(net898));
 sky130_fd_sc_hd__buf_8 fanout899 (.A(net900),
    .X(net899));
 sky130_fd_sc_hd__buf_8 fanout900 (.A(\ApproximateM_inst.lob_16.lob1.genblk1[2].genblk1.mux.sel ),
    .X(net900));
 sky130_fd_sc_hd__buf_8 fanout901 (.A(net902),
    .X(net901));
 sky130_fd_sc_hd__buf_12 fanout902 (.A(\ApproximateM_inst.lob_16.lob1.genblk1[1].genblk1.mux.sel ),
    .X(net902));
 sky130_fd_sc_hd__buf_4 fanout903 (.A(net904),
    .X(net903));
 sky130_fd_sc_hd__buf_8 fanout904 (.A(net909),
    .X(net904));
 sky130_fd_sc_hd__buf_4 fanout905 (.A(net906),
    .X(net905));
 sky130_fd_sc_hd__buf_2 fanout906 (.A(net909),
    .X(net906));
 sky130_fd_sc_hd__buf_4 fanout907 (.A(net908),
    .X(net907));
 sky130_fd_sc_hd__buf_6 fanout908 (.A(net909),
    .X(net908));
 sky130_fd_sc_hd__buf_4 fanout909 (.A(\ApproximateM_inst.lob_16.lob1.genblk1[1].genblk1.mux.sel ),
    .X(net909));
 sky130_fd_sc_hd__buf_8 fanout910 (.A(net912),
    .X(net910));
 sky130_fd_sc_hd__buf_4 fanout911 (.A(net912),
    .X(net911));
 sky130_fd_sc_hd__buf_8 fanout912 (.A(\ApproximateM_inst.lob_16.lob1.mux.sel ),
    .X(net912));
 sky130_fd_sc_hd__buf_8 fanout913 (.A(net918),
    .X(net913));
 sky130_fd_sc_hd__buf_4 fanout914 (.A(net915),
    .X(net914));
 sky130_fd_sc_hd__buf_4 fanout915 (.A(net917),
    .X(net915));
 sky130_fd_sc_hd__clkbuf_16 fanout916 (.A(net917),
    .X(net916));
 sky130_fd_sc_hd__clkbuf_4 fanout917 (.A(net918),
    .X(net917));
 sky130_fd_sc_hd__buf_6 fanout918 (.A(\ApproximateM_inst.lob_16.lob1.mux.sel ),
    .X(net918));
 sky130_fd_sc_hd__buf_6 fanout919 (.A(net922),
    .X(net919));
 sky130_fd_sc_hd__buf_4 fanout920 (.A(net921),
    .X(net920));
 sky130_fd_sc_hd__buf_4 fanout921 (.A(net922),
    .X(net921));
 sky130_fd_sc_hd__buf_4 fanout922 (.A(_08378_),
    .X(net922));
 sky130_fd_sc_hd__clkbuf_8 fanout923 (.A(net926),
    .X(net923));
 sky130_fd_sc_hd__buf_4 fanout924 (.A(net925),
    .X(net924));
 sky130_fd_sc_hd__clkbuf_8 fanout925 (.A(net926),
    .X(net925));
 sky130_fd_sc_hd__buf_4 fanout926 (.A(_08377_),
    .X(net926));
 sky130_fd_sc_hd__buf_4 fanout927 (.A(net930),
    .X(net927));
 sky130_fd_sc_hd__buf_2 fanout928 (.A(net930),
    .X(net928));
 sky130_fd_sc_hd__buf_4 fanout929 (.A(net930),
    .X(net929));
 sky130_fd_sc_hd__buf_2 fanout930 (.A(net935),
    .X(net930));
 sky130_fd_sc_hd__buf_4 fanout931 (.A(net932),
    .X(net931));
 sky130_fd_sc_hd__buf_4 fanout932 (.A(net935),
    .X(net932));
 sky130_fd_sc_hd__buf_4 fanout933 (.A(net934),
    .X(net933));
 sky130_fd_sc_hd__buf_4 fanout934 (.A(net935),
    .X(net934));
 sky130_fd_sc_hd__buf_4 fanout935 (.A(_03324_),
    .X(net935));
 sky130_fd_sc_hd__buf_4 fanout936 (.A(net937),
    .X(net936));
 sky130_fd_sc_hd__buf_4 fanout937 (.A(net938),
    .X(net937));
 sky130_fd_sc_hd__clkbuf_4 fanout938 (.A(_03324_),
    .X(net938));
 sky130_fd_sc_hd__buf_4 input1 (.A(buttons),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(i_wb_addr[17]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(i_wb_addr[18]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(i_wb_addr[19]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input13 (.A(i_wb_addr[1]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(i_wb_addr[20]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(i_wb_addr[21]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(i_wb_addr[22]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(i_wb_addr[23]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(i_wb_addr[24]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(i_wb_addr[25]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input2 (.A(i_wb_addr[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(i_wb_addr[26]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(i_wb_addr[27]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(i_wb_addr[28]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(i_wb_addr[29]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_8 input24 (.A(i_wb_addr[2]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(i_wb_addr[30]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(i_wb_addr[31]),
    .X(net26));
 sky130_fd_sc_hd__buf_6 input27 (.A(i_wb_addr[3]),
    .X(net27));
 sky130_fd_sc_hd__buf_4 input28 (.A(i_wb_addr[4]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(i_wb_addr[5]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(i_wb_addr[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(i_wb_addr[6]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(i_wb_addr[7]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(i_wb_addr[8]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(i_wb_addr[9]),
    .X(net33));
 sky130_fd_sc_hd__buf_8 input34 (.A(i_wb_cyc),
    .X(net34));
 sky130_fd_sc_hd__buf_4 input35 (.A(i_wb_data[0]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(i_wb_data[10]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(i_wb_data[11]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(i_wb_data[12]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(i_wb_data[13]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(i_wb_addr[11]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(i_wb_data[14]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(i_wb_data[15]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(i_wb_data[16]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(i_wb_data[17]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(i_wb_data[18]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(i_wb_data[19]),
    .X(net45));
 sky130_fd_sc_hd__buf_4 input46 (.A(i_wb_data[1]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(i_wb_data[20]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(i_wb_data[21]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(i_wb_data[22]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(i_wb_addr[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(i_wb_data[23]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(i_wb_data[24]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(i_wb_data[25]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(i_wb_data[26]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(i_wb_data[27]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(i_wb_data[28]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(i_wb_data[29]),
    .X(net56));
 sky130_fd_sc_hd__buf_4 input57 (.A(i_wb_data[2]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(i_wb_data[30]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(i_wb_data[31]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(i_wb_addr[13]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input60 (.A(i_wb_data[3]),
    .X(net60));
 sky130_fd_sc_hd__buf_2 input61 (.A(i_wb_data[4]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(i_wb_data[5]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 input63 (.A(i_wb_data[6]),
    .X(net63));
 sky130_fd_sc_hd__buf_2 input64 (.A(i_wb_data[7]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(i_wb_data[8]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 input66 (.A(i_wb_data[9]),
    .X(net66));
 sky130_fd_sc_hd__buf_8 input67 (.A(i_wb_stb),
    .X(net67));
 sky130_fd_sc_hd__buf_6 input68 (.A(i_wb_we),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_4 input69 (.A(reset),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(i_wb_addr[14]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(i_wb_addr[15]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(i_wb_addr[16]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 max_cap117 (.A(_04621_),
    .X(net117));
 sky130_fd_sc_hd__buf_2 max_cap118 (.A(_00184_),
    .X(net118));
 sky130_fd_sc_hd__buf_4 max_cap119 (.A(_02743_),
    .X(net119));
 sky130_fd_sc_hd__buf_4 max_cap121 (.A(_05241_),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_4 max_cap122 (.A(_01295_),
    .X(net122));
 sky130_fd_sc_hd__buf_6 max_cap139 (.A(_06098_),
    .X(net139));
 sky130_fd_sc_hd__buf_6 max_cap193 (.A(_06313_),
    .X(net193));
 sky130_fd_sc_hd__buf_6 max_cap197 (.A(_06245_),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 max_cap216 (.A(net217),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_2 max_cap217 (.A(_02595_),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_2 output100 (.A(net100),
    .X(o_wb_data[25]));
 sky130_fd_sc_hd__clkbuf_2 output101 (.A(net101),
    .X(o_wb_data[26]));
 sky130_fd_sc_hd__clkbuf_2 output102 (.A(net102),
    .X(o_wb_data[27]));
 sky130_fd_sc_hd__clkbuf_2 output103 (.A(net103),
    .X(o_wb_data[28]));
 sky130_fd_sc_hd__clkbuf_2 output104 (.A(net104),
    .X(o_wb_data[29]));
 sky130_fd_sc_hd__clkbuf_2 output105 (.A(net105),
    .X(o_wb_data[2]));
 sky130_fd_sc_hd__clkbuf_2 output106 (.A(net106),
    .X(o_wb_data[30]));
 sky130_fd_sc_hd__clkbuf_2 output107 (.A(net107),
    .X(o_wb_data[31]));
 sky130_fd_sc_hd__clkbuf_2 output108 (.A(net108),
    .X(o_wb_data[3]));
 sky130_fd_sc_hd__clkbuf_2 output109 (.A(net109),
    .X(o_wb_data[4]));
 sky130_fd_sc_hd__clkbuf_2 output110 (.A(net110),
    .X(o_wb_data[5]));
 sky130_fd_sc_hd__clkbuf_2 output111 (.A(net111),
    .X(o_wb_data[6]));
 sky130_fd_sc_hd__clkbuf_2 output112 (.A(net112),
    .X(o_wb_data[7]));
 sky130_fd_sc_hd__clkbuf_2 output113 (.A(net113),
    .X(o_wb_data[8]));
 sky130_fd_sc_hd__clkbuf_2 output114 (.A(net114),
    .X(o_wb_data[9]));
 sky130_fd_sc_hd__clkbuf_2 output70 (.A(net70),
    .X(leds[0]));
 sky130_fd_sc_hd__clkbuf_2 output71 (.A(net71),
    .X(leds[10]));
 sky130_fd_sc_hd__clkbuf_2 output72 (.A(net72),
    .X(leds[11]));
 sky130_fd_sc_hd__clkbuf_2 output73 (.A(net73),
    .X(leds[1]));
 sky130_fd_sc_hd__clkbuf_2 output74 (.A(net74),
    .X(leds[2]));
 sky130_fd_sc_hd__clkbuf_2 output75 (.A(net75),
    .X(leds[3]));
 sky130_fd_sc_hd__clkbuf_2 output76 (.A(net76),
    .X(leds[4]));
 sky130_fd_sc_hd__clkbuf_2 output77 (.A(net77),
    .X(leds[5]));
 sky130_fd_sc_hd__clkbuf_2 output78 (.A(net78),
    .X(leds[6]));
 sky130_fd_sc_hd__clkbuf_2 output79 (.A(net79),
    .X(leds[7]));
 sky130_fd_sc_hd__clkbuf_2 output80 (.A(net80),
    .X(leds[8]));
 sky130_fd_sc_hd__clkbuf_2 output81 (.A(net81),
    .X(leds[9]));
 sky130_fd_sc_hd__clkbuf_2 output82 (.A(net82),
    .X(o_wb_ack));
 sky130_fd_sc_hd__clkbuf_2 output83 (.A(net83),
    .X(o_wb_data[0]));
 sky130_fd_sc_hd__clkbuf_2 output84 (.A(net84),
    .X(o_wb_data[10]));
 sky130_fd_sc_hd__clkbuf_2 output85 (.A(net85),
    .X(o_wb_data[11]));
 sky130_fd_sc_hd__clkbuf_2 output86 (.A(net86),
    .X(o_wb_data[12]));
 sky130_fd_sc_hd__clkbuf_2 output87 (.A(net87),
    .X(o_wb_data[13]));
 sky130_fd_sc_hd__clkbuf_2 output88 (.A(net88),
    .X(o_wb_data[14]));
 sky130_fd_sc_hd__clkbuf_2 output89 (.A(net89),
    .X(o_wb_data[15]));
 sky130_fd_sc_hd__clkbuf_2 output90 (.A(net90),
    .X(o_wb_data[16]));
 sky130_fd_sc_hd__clkbuf_2 output91 (.A(net91),
    .X(o_wb_data[17]));
 sky130_fd_sc_hd__clkbuf_2 output92 (.A(net92),
    .X(o_wb_data[18]));
 sky130_fd_sc_hd__clkbuf_2 output93 (.A(net93),
    .X(o_wb_data[19]));
 sky130_fd_sc_hd__clkbuf_2 output94 (.A(net94),
    .X(o_wb_data[1]));
 sky130_fd_sc_hd__clkbuf_2 output95 (.A(net95),
    .X(o_wb_data[20]));
 sky130_fd_sc_hd__clkbuf_2 output96 (.A(net96),
    .X(o_wb_data[21]));
 sky130_fd_sc_hd__clkbuf_2 output97 (.A(net97),
    .X(o_wb_data[22]));
 sky130_fd_sc_hd__clkbuf_2 output98 (.A(net98),
    .X(o_wb_data[23]));
 sky130_fd_sc_hd__clkbuf_2 output99 (.A(net99),
    .X(o_wb_data[24]));
 sky130_fd_sc_hd__conb_1 wb_buttons_leds_939 (.LO(net939));
 sky130_fd_sc_hd__conb_1 wb_buttons_leds_940 (.LO(net940));
 sky130_fd_sc_hd__conb_1 wb_buttons_leds_941 (.LO(net941));
 sky130_fd_sc_hd__conb_1 wb_buttons_leds_942 (.LO(net942));
 sky130_fd_sc_hd__conb_1 wb_buttons_leds_943 (.LO(net943));
 sky130_fd_sc_hd__conb_1 wb_buttons_leds_944 (.LO(net944));
 sky130_fd_sc_hd__conb_1 wb_buttons_leds_945 (.LO(net945));
 sky130_fd_sc_hd__conb_1 wb_buttons_leds_946 (.LO(net946));
 sky130_fd_sc_hd__conb_1 wb_buttons_leds_947 (.LO(net947));
 sky130_fd_sc_hd__conb_1 wb_buttons_leds_948 (.LO(net948));
 sky130_fd_sc_hd__conb_1 wb_buttons_leds_949 (.LO(net949));
 sky130_fd_sc_hd__conb_1 wb_buttons_leds_950 (.LO(net950));
 sky130_fd_sc_hd__conb_1 wb_buttons_leds_951 (.LO(net951));
 sky130_fd_sc_hd__buf_2 wire115 (.A(_04869_),
    .X(net115));
 sky130_fd_sc_hd__buf_4 wire116 (.A(_03343_),
    .X(net116));
 sky130_fd_sc_hd__buf_4 wire120 (.A(_01428_),
    .X(net120));
 sky130_fd_sc_hd__buf_2 wire222 (.A(_08388_),
    .X(net222));
 sky130_fd_sc_hd__buf_4 wire268 (.A(_06169_),
    .X(net268));
 assign led_enb[0] = net939;
 assign led_enb[10] = net949;
 assign led_enb[11] = net950;
 assign led_enb[1] = net940;
 assign led_enb[2] = net941;
 assign led_enb[3] = net942;
 assign led_enb[4] = net943;
 assign led_enb[5] = net944;
 assign led_enb[6] = net945;
 assign led_enb[7] = net946;
 assign led_enb[8] = net947;
 assign led_enb[9] = net948;
 assign o_wb_stall = net951;
endmodule

