magic
tech sky130A
magscale 1 2
timestamp 1698766093
<< obsli1 >>
rect 1104 2159 108836 107729
<< obsm1 >>
rect 934 892 109098 107760
<< metal2 >>
rect 27434 109200 27490 110000
rect 82450 109200 82506 110000
rect 3054 0 3110 800
rect 7378 0 7434 800
rect 11702 0 11758 800
rect 16026 0 16082 800
rect 20350 0 20406 800
rect 24674 0 24730 800
rect 28998 0 29054 800
rect 33322 0 33378 800
rect 37646 0 37702 800
rect 41970 0 42026 800
rect 46294 0 46350 800
rect 50618 0 50674 800
rect 54942 0 54998 800
rect 59266 0 59322 800
rect 63590 0 63646 800
rect 67914 0 67970 800
rect 72238 0 72294 800
rect 76562 0 76618 800
rect 80886 0 80942 800
rect 85210 0 85266 800
rect 89534 0 89590 800
rect 93858 0 93914 800
rect 98182 0 98238 800
rect 102506 0 102562 800
rect 106830 0 106886 800
<< obsm2 >>
rect 938 109144 27378 109200
rect 27546 109144 82394 109200
rect 82562 109144 109094 109200
rect 938 856 109094 109144
rect 938 800 2998 856
rect 3166 800 7322 856
rect 7490 800 11646 856
rect 11814 800 15970 856
rect 16138 800 20294 856
rect 20462 800 24618 856
rect 24786 800 28942 856
rect 29110 800 33266 856
rect 33434 800 37590 856
rect 37758 800 41914 856
rect 42082 800 46238 856
rect 46406 800 50562 856
rect 50730 800 54886 856
rect 55054 800 59210 856
rect 59378 800 63534 856
rect 63702 800 67858 856
rect 68026 800 72182 856
rect 72350 800 76506 856
rect 76674 800 80830 856
rect 80998 800 85154 856
rect 85322 800 89478 856
rect 89646 800 93802 856
rect 93970 800 98126 856
rect 98294 800 102450 856
rect 102618 800 106774 856
rect 106942 800 109094 856
<< metal3 >>
rect 0 106632 800 106752
rect 0 105544 800 105664
rect 0 104456 800 104576
rect 0 103368 800 103488
rect 0 102280 800 102400
rect 0 101192 800 101312
rect 0 100104 800 100224
rect 0 99016 800 99136
rect 109200 98744 110000 98864
rect 0 97928 800 98048
rect 0 96840 800 96960
rect 0 95752 800 95872
rect 0 94664 800 94784
rect 0 93576 800 93696
rect 0 92488 800 92608
rect 0 91400 800 91520
rect 0 90312 800 90432
rect 0 89224 800 89344
rect 0 88136 800 88256
rect 0 87048 800 87168
rect 0 85960 800 86080
rect 0 84872 800 84992
rect 0 83784 800 83904
rect 0 82696 800 82816
rect 0 81608 800 81728
rect 0 80520 800 80640
rect 0 79432 800 79552
rect 0 78344 800 78464
rect 0 77256 800 77376
rect 109200 76848 110000 76968
rect 0 76168 800 76288
rect 0 75080 800 75200
rect 0 73992 800 74112
rect 0 72904 800 73024
rect 0 71816 800 71936
rect 0 70728 800 70848
rect 0 69640 800 69760
rect 0 68552 800 68672
rect 0 67464 800 67584
rect 0 66376 800 66496
rect 0 65288 800 65408
rect 0 64200 800 64320
rect 0 63112 800 63232
rect 0 62024 800 62144
rect 0 60936 800 61056
rect 0 59848 800 59968
rect 0 58760 800 58880
rect 0 57672 800 57792
rect 0 56584 800 56704
rect 0 55496 800 55616
rect 109200 54952 110000 55072
rect 0 54408 800 54528
rect 0 53320 800 53440
rect 0 52232 800 52352
rect 0 51144 800 51264
rect 0 50056 800 50176
rect 0 48968 800 49088
rect 0 47880 800 48000
rect 0 46792 800 46912
rect 0 45704 800 45824
rect 0 44616 800 44736
rect 0 43528 800 43648
rect 0 42440 800 42560
rect 0 41352 800 41472
rect 0 40264 800 40384
rect 0 39176 800 39296
rect 0 38088 800 38208
rect 0 37000 800 37120
rect 0 35912 800 36032
rect 0 34824 800 34944
rect 0 33736 800 33856
rect 109200 33056 110000 33176
rect 0 32648 800 32768
rect 0 31560 800 31680
rect 0 30472 800 30592
rect 0 29384 800 29504
rect 0 28296 800 28416
rect 0 27208 800 27328
rect 0 26120 800 26240
rect 0 25032 800 25152
rect 0 23944 800 24064
rect 0 22856 800 22976
rect 0 21768 800 21888
rect 0 20680 800 20800
rect 0 19592 800 19712
rect 0 18504 800 18624
rect 0 17416 800 17536
rect 0 16328 800 16448
rect 0 15240 800 15360
rect 0 14152 800 14272
rect 0 13064 800 13184
rect 0 11976 800 12096
rect 109200 11160 110000 11280
rect 0 10888 800 11008
rect 0 9800 800 9920
rect 0 8712 800 8832
rect 0 7624 800 7744
rect 0 6536 800 6656
rect 0 5448 800 5568
rect 0 4360 800 4480
rect 0 3272 800 3392
<< obsm3 >>
rect 800 106832 109200 107745
rect 880 106552 109200 106832
rect 800 105744 109200 106552
rect 880 105464 109200 105744
rect 800 104656 109200 105464
rect 880 104376 109200 104656
rect 800 103568 109200 104376
rect 880 103288 109200 103568
rect 800 102480 109200 103288
rect 880 102200 109200 102480
rect 800 101392 109200 102200
rect 880 101112 109200 101392
rect 800 100304 109200 101112
rect 880 100024 109200 100304
rect 800 99216 109200 100024
rect 880 98944 109200 99216
rect 880 98936 109120 98944
rect 800 98664 109120 98936
rect 800 98128 109200 98664
rect 880 97848 109200 98128
rect 800 97040 109200 97848
rect 880 96760 109200 97040
rect 800 95952 109200 96760
rect 880 95672 109200 95952
rect 800 94864 109200 95672
rect 880 94584 109200 94864
rect 800 93776 109200 94584
rect 880 93496 109200 93776
rect 800 92688 109200 93496
rect 880 92408 109200 92688
rect 800 91600 109200 92408
rect 880 91320 109200 91600
rect 800 90512 109200 91320
rect 880 90232 109200 90512
rect 800 89424 109200 90232
rect 880 89144 109200 89424
rect 800 88336 109200 89144
rect 880 88056 109200 88336
rect 800 87248 109200 88056
rect 880 86968 109200 87248
rect 800 86160 109200 86968
rect 880 85880 109200 86160
rect 800 85072 109200 85880
rect 880 84792 109200 85072
rect 800 83984 109200 84792
rect 880 83704 109200 83984
rect 800 82896 109200 83704
rect 880 82616 109200 82896
rect 800 81808 109200 82616
rect 880 81528 109200 81808
rect 800 80720 109200 81528
rect 880 80440 109200 80720
rect 800 79632 109200 80440
rect 880 79352 109200 79632
rect 800 78544 109200 79352
rect 880 78264 109200 78544
rect 800 77456 109200 78264
rect 880 77176 109200 77456
rect 800 77048 109200 77176
rect 800 76768 109120 77048
rect 800 76368 109200 76768
rect 880 76088 109200 76368
rect 800 75280 109200 76088
rect 880 75000 109200 75280
rect 800 74192 109200 75000
rect 880 73912 109200 74192
rect 800 73104 109200 73912
rect 880 72824 109200 73104
rect 800 72016 109200 72824
rect 880 71736 109200 72016
rect 800 70928 109200 71736
rect 880 70648 109200 70928
rect 800 69840 109200 70648
rect 880 69560 109200 69840
rect 800 68752 109200 69560
rect 880 68472 109200 68752
rect 800 67664 109200 68472
rect 880 67384 109200 67664
rect 800 66576 109200 67384
rect 880 66296 109200 66576
rect 800 65488 109200 66296
rect 880 65208 109200 65488
rect 800 64400 109200 65208
rect 880 64120 109200 64400
rect 800 63312 109200 64120
rect 880 63032 109200 63312
rect 800 62224 109200 63032
rect 880 61944 109200 62224
rect 800 61136 109200 61944
rect 880 60856 109200 61136
rect 800 60048 109200 60856
rect 880 59768 109200 60048
rect 800 58960 109200 59768
rect 880 58680 109200 58960
rect 800 57872 109200 58680
rect 880 57592 109200 57872
rect 800 56784 109200 57592
rect 880 56504 109200 56784
rect 800 55696 109200 56504
rect 880 55416 109200 55696
rect 800 55152 109200 55416
rect 800 54872 109120 55152
rect 800 54608 109200 54872
rect 880 54328 109200 54608
rect 800 53520 109200 54328
rect 880 53240 109200 53520
rect 800 52432 109200 53240
rect 880 52152 109200 52432
rect 800 51344 109200 52152
rect 880 51064 109200 51344
rect 800 50256 109200 51064
rect 880 49976 109200 50256
rect 800 49168 109200 49976
rect 880 48888 109200 49168
rect 800 48080 109200 48888
rect 880 47800 109200 48080
rect 800 46992 109200 47800
rect 880 46712 109200 46992
rect 800 45904 109200 46712
rect 880 45624 109200 45904
rect 800 44816 109200 45624
rect 880 44536 109200 44816
rect 800 43728 109200 44536
rect 880 43448 109200 43728
rect 800 42640 109200 43448
rect 880 42360 109200 42640
rect 800 41552 109200 42360
rect 880 41272 109200 41552
rect 800 40464 109200 41272
rect 880 40184 109200 40464
rect 800 39376 109200 40184
rect 880 39096 109200 39376
rect 800 38288 109200 39096
rect 880 38008 109200 38288
rect 800 37200 109200 38008
rect 880 36920 109200 37200
rect 800 36112 109200 36920
rect 880 35832 109200 36112
rect 800 35024 109200 35832
rect 880 34744 109200 35024
rect 800 33936 109200 34744
rect 880 33656 109200 33936
rect 800 33256 109200 33656
rect 800 32976 109120 33256
rect 800 32848 109200 32976
rect 880 32568 109200 32848
rect 800 31760 109200 32568
rect 880 31480 109200 31760
rect 800 30672 109200 31480
rect 880 30392 109200 30672
rect 800 29584 109200 30392
rect 880 29304 109200 29584
rect 800 28496 109200 29304
rect 880 28216 109200 28496
rect 800 27408 109200 28216
rect 880 27128 109200 27408
rect 800 26320 109200 27128
rect 880 26040 109200 26320
rect 800 25232 109200 26040
rect 880 24952 109200 25232
rect 800 24144 109200 24952
rect 880 23864 109200 24144
rect 800 23056 109200 23864
rect 880 22776 109200 23056
rect 800 21968 109200 22776
rect 880 21688 109200 21968
rect 800 20880 109200 21688
rect 880 20600 109200 20880
rect 800 19792 109200 20600
rect 880 19512 109200 19792
rect 800 18704 109200 19512
rect 880 18424 109200 18704
rect 800 17616 109200 18424
rect 880 17336 109200 17616
rect 800 16528 109200 17336
rect 880 16248 109200 16528
rect 800 15440 109200 16248
rect 880 15160 109200 15440
rect 800 14352 109200 15160
rect 880 14072 109200 14352
rect 800 13264 109200 14072
rect 880 12984 109200 13264
rect 800 12176 109200 12984
rect 880 11896 109200 12176
rect 800 11360 109200 11896
rect 800 11088 109120 11360
rect 880 11080 109120 11088
rect 880 10808 109200 11080
rect 800 10000 109200 10808
rect 880 9720 109200 10000
rect 800 8912 109200 9720
rect 880 8632 109200 8912
rect 800 7824 109200 8632
rect 880 7544 109200 7824
rect 800 6736 109200 7544
rect 880 6456 109200 6736
rect 800 5648 109200 6456
rect 880 5368 109200 5648
rect 800 4560 109200 5368
rect 880 4280 109200 4560
rect 800 3472 109200 4280
rect 880 3192 109200 3472
rect 800 2143 109200 3192
<< metal4 >>
rect 4208 2128 4528 107760
rect 19568 2128 19888 107760
rect 34928 2128 35248 107760
rect 50288 2128 50608 107760
rect 65648 2128 65968 107760
rect 81008 2128 81328 107760
rect 96368 2128 96688 107760
<< obsm4 >>
rect 3003 2347 4128 106317
rect 4608 2347 19488 106317
rect 19968 2347 34848 106317
rect 35328 2347 50208 106317
rect 50688 2347 65568 106317
rect 66048 2347 80928 106317
rect 81408 2347 93965 106317
<< labels >>
rlabel metal2 s 3054 0 3110 800 6 buttons
port 1 nsew signal input
rlabel metal2 s 82450 109200 82506 110000 6 clk
port 2 nsew signal input
rlabel metal3 s 0 3272 800 3392 6 i_wb_addr[0]
port 3 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 i_wb_addr[10]
port 4 nsew signal input
rlabel metal3 s 0 15240 800 15360 6 i_wb_addr[11]
port 5 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 i_wb_addr[12]
port 6 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 i_wb_addr[13]
port 7 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 i_wb_addr[14]
port 8 nsew signal input
rlabel metal3 s 0 19592 800 19712 6 i_wb_addr[15]
port 9 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 i_wb_addr[16]
port 10 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 i_wb_addr[17]
port 11 nsew signal input
rlabel metal3 s 0 22856 800 22976 6 i_wb_addr[18]
port 12 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 i_wb_addr[19]
port 13 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 i_wb_addr[1]
port 14 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 i_wb_addr[20]
port 15 nsew signal input
rlabel metal3 s 0 26120 800 26240 6 i_wb_addr[21]
port 16 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 i_wb_addr[22]
port 17 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 i_wb_addr[23]
port 18 nsew signal input
rlabel metal3 s 0 29384 800 29504 6 i_wb_addr[24]
port 19 nsew signal input
rlabel metal3 s 0 30472 800 30592 6 i_wb_addr[25]
port 20 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 i_wb_addr[26]
port 21 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 i_wb_addr[27]
port 22 nsew signal input
rlabel metal3 s 0 33736 800 33856 6 i_wb_addr[28]
port 23 nsew signal input
rlabel metal3 s 0 34824 800 34944 6 i_wb_addr[29]
port 24 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 i_wb_addr[2]
port 25 nsew signal input
rlabel metal3 s 0 35912 800 36032 6 i_wb_addr[30]
port 26 nsew signal input
rlabel metal3 s 0 37000 800 37120 6 i_wb_addr[31]
port 27 nsew signal input
rlabel metal3 s 0 6536 800 6656 6 i_wb_addr[3]
port 28 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 i_wb_addr[4]
port 29 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 i_wb_addr[5]
port 30 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 i_wb_addr[6]
port 31 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 i_wb_addr[7]
port 32 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 i_wb_addr[8]
port 33 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 i_wb_addr[9]
port 34 nsew signal input
rlabel metal3 s 109200 11160 110000 11280 6 i_wb_cyc
port 35 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 i_wb_data[0]
port 36 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 i_wb_data[10]
port 37 nsew signal input
rlabel metal3 s 0 50056 800 50176 6 i_wb_data[11]
port 38 nsew signal input
rlabel metal3 s 0 51144 800 51264 6 i_wb_data[12]
port 39 nsew signal input
rlabel metal3 s 0 52232 800 52352 6 i_wb_data[13]
port 40 nsew signal input
rlabel metal3 s 0 53320 800 53440 6 i_wb_data[14]
port 41 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 i_wb_data[15]
port 42 nsew signal input
rlabel metal3 s 0 55496 800 55616 6 i_wb_data[16]
port 43 nsew signal input
rlabel metal3 s 0 56584 800 56704 6 i_wb_data[17]
port 44 nsew signal input
rlabel metal3 s 0 57672 800 57792 6 i_wb_data[18]
port 45 nsew signal input
rlabel metal3 s 0 58760 800 58880 6 i_wb_data[19]
port 46 nsew signal input
rlabel metal3 s 0 39176 800 39296 6 i_wb_data[1]
port 47 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 i_wb_data[20]
port 48 nsew signal input
rlabel metal3 s 0 60936 800 61056 6 i_wb_data[21]
port 49 nsew signal input
rlabel metal3 s 0 62024 800 62144 6 i_wb_data[22]
port 50 nsew signal input
rlabel metal3 s 0 63112 800 63232 6 i_wb_data[23]
port 51 nsew signal input
rlabel metal3 s 0 64200 800 64320 6 i_wb_data[24]
port 52 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 i_wb_data[25]
port 53 nsew signal input
rlabel metal3 s 0 66376 800 66496 6 i_wb_data[26]
port 54 nsew signal input
rlabel metal3 s 0 67464 800 67584 6 i_wb_data[27]
port 55 nsew signal input
rlabel metal3 s 0 68552 800 68672 6 i_wb_data[28]
port 56 nsew signal input
rlabel metal3 s 0 69640 800 69760 6 i_wb_data[29]
port 57 nsew signal input
rlabel metal3 s 0 40264 800 40384 6 i_wb_data[2]
port 58 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 i_wb_data[30]
port 59 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 i_wb_data[31]
port 60 nsew signal input
rlabel metal3 s 0 41352 800 41472 6 i_wb_data[3]
port 61 nsew signal input
rlabel metal3 s 0 42440 800 42560 6 i_wb_data[4]
port 62 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 i_wb_data[5]
port 63 nsew signal input
rlabel metal3 s 0 44616 800 44736 6 i_wb_data[6]
port 64 nsew signal input
rlabel metal3 s 0 45704 800 45824 6 i_wb_data[7]
port 65 nsew signal input
rlabel metal3 s 0 46792 800 46912 6 i_wb_data[8]
port 66 nsew signal input
rlabel metal3 s 0 47880 800 48000 6 i_wb_data[9]
port 67 nsew signal input
rlabel metal3 s 109200 33056 110000 33176 6 i_wb_stb
port 68 nsew signal input
rlabel metal3 s 109200 54952 110000 55072 6 i_wb_we
port 69 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 led_enb[0]
port 70 nsew signal output
rlabel metal2 s 50618 0 50674 800 6 led_enb[10]
port 71 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 led_enb[11]
port 72 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 led_enb[1]
port 73 nsew signal output
rlabel metal2 s 16026 0 16082 800 6 led_enb[2]
port 74 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 led_enb[3]
port 75 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 led_enb[4]
port 76 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 led_enb[5]
port 77 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 led_enb[6]
port 78 nsew signal output
rlabel metal2 s 37646 0 37702 800 6 led_enb[7]
port 79 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 led_enb[8]
port 80 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 led_enb[9]
port 81 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 leds[0]
port 82 nsew signal output
rlabel metal2 s 102506 0 102562 800 6 leds[10]
port 83 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 leds[11]
port 84 nsew signal output
rlabel metal2 s 63590 0 63646 800 6 leds[1]
port 85 nsew signal output
rlabel metal2 s 67914 0 67970 800 6 leds[2]
port 86 nsew signal output
rlabel metal2 s 72238 0 72294 800 6 leds[3]
port 87 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 leds[4]
port 88 nsew signal output
rlabel metal2 s 80886 0 80942 800 6 leds[5]
port 89 nsew signal output
rlabel metal2 s 85210 0 85266 800 6 leds[6]
port 90 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 leds[7]
port 91 nsew signal output
rlabel metal2 s 93858 0 93914 800 6 leds[8]
port 92 nsew signal output
rlabel metal2 s 98182 0 98238 800 6 leds[9]
port 93 nsew signal output
rlabel metal3 s 109200 76848 110000 76968 6 o_wb_ack
port 94 nsew signal output
rlabel metal3 s 0 72904 800 73024 6 o_wb_data[0]
port 95 nsew signal output
rlabel metal3 s 0 83784 800 83904 6 o_wb_data[10]
port 96 nsew signal output
rlabel metal3 s 0 84872 800 84992 6 o_wb_data[11]
port 97 nsew signal output
rlabel metal3 s 0 85960 800 86080 6 o_wb_data[12]
port 98 nsew signal output
rlabel metal3 s 0 87048 800 87168 6 o_wb_data[13]
port 99 nsew signal output
rlabel metal3 s 0 88136 800 88256 6 o_wb_data[14]
port 100 nsew signal output
rlabel metal3 s 0 89224 800 89344 6 o_wb_data[15]
port 101 nsew signal output
rlabel metal3 s 0 90312 800 90432 6 o_wb_data[16]
port 102 nsew signal output
rlabel metal3 s 0 91400 800 91520 6 o_wb_data[17]
port 103 nsew signal output
rlabel metal3 s 0 92488 800 92608 6 o_wb_data[18]
port 104 nsew signal output
rlabel metal3 s 0 93576 800 93696 6 o_wb_data[19]
port 105 nsew signal output
rlabel metal3 s 0 73992 800 74112 6 o_wb_data[1]
port 106 nsew signal output
rlabel metal3 s 0 94664 800 94784 6 o_wb_data[20]
port 107 nsew signal output
rlabel metal3 s 0 95752 800 95872 6 o_wb_data[21]
port 108 nsew signal output
rlabel metal3 s 0 96840 800 96960 6 o_wb_data[22]
port 109 nsew signal output
rlabel metal3 s 0 97928 800 98048 6 o_wb_data[23]
port 110 nsew signal output
rlabel metal3 s 0 99016 800 99136 6 o_wb_data[24]
port 111 nsew signal output
rlabel metal3 s 0 100104 800 100224 6 o_wb_data[25]
port 112 nsew signal output
rlabel metal3 s 0 101192 800 101312 6 o_wb_data[26]
port 113 nsew signal output
rlabel metal3 s 0 102280 800 102400 6 o_wb_data[27]
port 114 nsew signal output
rlabel metal3 s 0 103368 800 103488 6 o_wb_data[28]
port 115 nsew signal output
rlabel metal3 s 0 104456 800 104576 6 o_wb_data[29]
port 116 nsew signal output
rlabel metal3 s 0 75080 800 75200 6 o_wb_data[2]
port 117 nsew signal output
rlabel metal3 s 0 105544 800 105664 6 o_wb_data[30]
port 118 nsew signal output
rlabel metal3 s 0 106632 800 106752 6 o_wb_data[31]
port 119 nsew signal output
rlabel metal3 s 0 76168 800 76288 6 o_wb_data[3]
port 120 nsew signal output
rlabel metal3 s 0 77256 800 77376 6 o_wb_data[4]
port 121 nsew signal output
rlabel metal3 s 0 78344 800 78464 6 o_wb_data[5]
port 122 nsew signal output
rlabel metal3 s 0 79432 800 79552 6 o_wb_data[6]
port 123 nsew signal output
rlabel metal3 s 0 80520 800 80640 6 o_wb_data[7]
port 124 nsew signal output
rlabel metal3 s 0 81608 800 81728 6 o_wb_data[8]
port 125 nsew signal output
rlabel metal3 s 0 82696 800 82816 6 o_wb_data[9]
port 126 nsew signal output
rlabel metal3 s 109200 98744 110000 98864 6 o_wb_stall
port 127 nsew signal output
rlabel metal2 s 27434 109200 27490 110000 6 reset
port 128 nsew signal input
rlabel metal4 s 4208 2128 4528 107760 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 107760 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 107760 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 107760 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 107760 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 107760 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 107760 6 vssd1
port 130 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 110000 110000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 27395712
string GDS_FILE /home/bignixon/unic-cass/caravel_tutorial/caravel_user_project/openlane/wb_buttons_leds/runs/23_10_31_12_19/results/signoff/wb_buttons_leds.magic.gds
string GDS_START 1498246
<< end >>

