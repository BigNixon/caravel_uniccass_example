magic
tech sky130A
magscale 1 2
timestamp 1698268990
<< checkpaint >>
rect -12658 -11586 596582 715522
<< metal1 >>
rect 59170 2864 59176 2916
rect 59228 2904 59234 2916
rect 64552 2904 64558 2916
rect 59228 2876 64558 2904
rect 59228 2864 59234 2876
rect 64552 2864 64558 2876
rect 64610 2864 64616 2916
rect 67634 2864 67640 2916
rect 67692 2904 67698 2916
rect 70072 2904 70078 2916
rect 67692 2876 70078 2904
rect 67692 2864 67698 2876
rect 70072 2864 70078 2876
rect 70130 2864 70136 2916
rect 71774 2864 71780 2916
rect 71832 2904 71838 2916
rect 74488 2904 74494 2916
rect 71832 2876 74494 2904
rect 71832 2864 71838 2876
rect 74488 2864 74494 2876
rect 74546 2864 74552 2916
rect 75454 2864 75460 2916
rect 75512 2904 75518 2916
rect 76696 2904 76702 2916
rect 75512 2876 76702 2904
rect 75512 2864 75518 2876
rect 76696 2864 76702 2876
rect 76754 2864 76760 2916
rect 80146 2864 80152 2916
rect 80204 2904 80210 2916
rect 84424 2904 84430 2916
rect 80204 2876 84430 2904
rect 80204 2864 80210 2876
rect 84424 2864 84430 2876
rect 84482 2864 84488 2916
rect 85390 2864 85396 2916
rect 85448 2904 85454 2916
rect 86632 2904 86638 2916
rect 85448 2876 86638 2904
rect 85448 2864 85454 2876
rect 86632 2864 86638 2876
rect 86690 2864 86696 2916
rect 86770 2864 86776 2916
rect 86828 2904 86834 2916
rect 87736 2904 87742 2916
rect 86828 2876 87742 2904
rect 86828 2864 86834 2876
rect 87736 2864 87742 2876
rect 87794 2864 87800 2916
rect 88150 2864 88156 2916
rect 88208 2904 88214 2916
rect 92152 2904 92158 2916
rect 88208 2876 92158 2904
rect 88208 2864 88214 2876
rect 92152 2864 92158 2876
rect 92210 2864 92216 2916
rect 92474 2864 92480 2916
rect 92532 2904 92538 2916
rect 94360 2904 94366 2916
rect 92532 2876 94366 2904
rect 92532 2864 92538 2876
rect 94360 2864 94366 2876
rect 94418 2864 94424 2916
rect 94590 2864 94596 2916
rect 94648 2904 94654 2916
rect 95464 2904 95470 2916
rect 94648 2876 95470 2904
rect 94648 2864 94654 2876
rect 95464 2864 95470 2876
rect 95522 2864 95528 2916
rect 95694 2864 95700 2916
rect 95752 2904 95758 2916
rect 97672 2904 97678 2916
rect 95752 2876 97678 2904
rect 95752 2864 95758 2876
rect 97672 2864 97678 2876
rect 97730 2864 97736 2916
rect 97994 2864 98000 2916
rect 98052 2904 98058 2916
rect 100984 2904 100990 2916
rect 98052 2876 100990 2904
rect 98052 2864 98058 2876
rect 100984 2864 100990 2876
rect 101042 2864 101048 2916
rect 102226 2864 102232 2916
rect 102284 2904 102290 2916
rect 105400 2904 105406 2916
rect 102284 2876 105406 2904
rect 102284 2864 102290 2876
rect 105400 2864 105406 2876
rect 105458 2864 105464 2916
rect 105538 2864 105544 2916
rect 105596 2904 105602 2916
rect 106504 2904 106510 2916
rect 105596 2876 106510 2904
rect 105596 2864 105602 2876
rect 106504 2864 106510 2876
rect 106562 2864 106568 2916
rect 107746 2864 107752 2916
rect 107804 2904 107810 2916
rect 109816 2904 109822 2916
rect 107804 2876 109822 2904
rect 107804 2864 107810 2876
rect 109816 2864 109822 2876
rect 109874 2864 109880 2916
rect 110414 2864 110420 2916
rect 110472 2904 110478 2916
rect 113128 2904 113134 2916
rect 110472 2876 113134 2904
rect 110472 2864 110478 2876
rect 113128 2864 113134 2876
rect 113186 2864 113192 2916
rect 114738 2864 114744 2916
rect 114796 2904 114802 2916
rect 116440 2904 116446 2916
rect 114796 2876 116446 2904
rect 114796 2864 114802 2876
rect 116440 2864 116446 2876
rect 116498 2864 116504 2916
rect 117314 2864 117320 2916
rect 117372 2904 117378 2916
rect 119752 2904 119758 2916
rect 117372 2876 119758 2904
rect 117372 2864 117378 2876
rect 119752 2864 119758 2876
rect 119810 2864 119816 2916
rect 120074 2864 120080 2916
rect 120132 2904 120138 2916
rect 124168 2904 124174 2916
rect 120132 2876 124174 2904
rect 120132 2864 120138 2876
rect 124168 2864 124174 2876
rect 124226 2864 124232 2916
rect 125134 2864 125140 2916
rect 125192 2904 125198 2916
rect 127480 2904 127486 2916
rect 125192 2876 127486 2904
rect 125192 2864 125198 2876
rect 127480 2864 127486 2876
rect 127538 2864 127544 2916
rect 127618 2864 127624 2916
rect 127676 2904 127682 2916
rect 129688 2904 129694 2916
rect 127676 2876 129694 2904
rect 127676 2864 127682 2876
rect 129688 2864 129694 2876
rect 129746 2864 129752 2916
rect 133230 2864 133236 2916
rect 133288 2904 133294 2916
rect 134104 2904 134110 2916
rect 133288 2876 134110 2904
rect 133288 2864 133294 2876
rect 134104 2864 134110 2876
rect 134162 2864 134168 2916
rect 136634 2864 136640 2916
rect 136692 2904 136698 2916
rect 139624 2904 139630 2916
rect 136692 2876 139630 2904
rect 136692 2864 136698 2876
rect 139624 2864 139630 2876
rect 139682 2864 139688 2916
rect 144178 2864 144184 2916
rect 144236 2904 144242 2916
rect 146248 2904 146254 2916
rect 144236 2876 146254 2904
rect 144236 2864 144242 2876
rect 146248 2864 146254 2876
rect 146306 2864 146312 2916
rect 149054 2864 149060 2916
rect 149112 2904 149118 2916
rect 151768 2904 151774 2916
rect 149112 2876 151774 2904
rect 149112 2864 149118 2876
rect 151768 2864 151774 2876
rect 151826 2864 151832 2916
rect 153378 2864 153384 2916
rect 153436 2904 153442 2916
rect 155080 2904 155086 2916
rect 153436 2876 155086 2904
rect 153436 2864 153442 2876
rect 155080 2864 155086 2876
rect 155138 2864 155144 2916
rect 155954 2864 155960 2916
rect 156012 2904 156018 2916
rect 158392 2904 158398 2916
rect 156012 2876 158398 2904
rect 156012 2864 156018 2876
rect 158392 2864 158398 2876
rect 158450 2864 158456 2916
rect 158714 2864 158720 2916
rect 158772 2904 158778 2916
rect 162808 2904 162814 2916
rect 158772 2876 162814 2904
rect 158772 2864 158778 2876
rect 162808 2864 162814 2876
rect 162866 2864 162872 2916
rect 166994 2864 167000 2916
rect 167052 2904 167058 2916
rect 169432 2904 169438 2916
rect 167052 2876 169438 2904
rect 167052 2864 167058 2876
rect 169432 2864 169438 2876
rect 169490 2864 169496 2916
rect 169570 2864 169576 2916
rect 169628 2904 169634 2916
rect 170536 2904 170542 2916
rect 169628 2876 170542 2904
rect 169628 2864 169634 2876
rect 170536 2864 170542 2876
rect 170594 2864 170600 2916
rect 172974 2864 172980 2916
rect 173032 2904 173038 2916
rect 174952 2904 174958 2916
rect 173032 2876 174958 2904
rect 173032 2864 173038 2876
rect 174952 2864 174958 2876
rect 175010 2864 175016 2916
rect 175274 2864 175280 2916
rect 175332 2904 175338 2916
rect 178264 2904 178270 2916
rect 175332 2876 178270 2904
rect 175332 2864 175338 2876
rect 178264 2864 178270 2876
rect 178322 2864 178328 2916
rect 179506 2864 179512 2916
rect 179564 2904 179570 2916
rect 181576 2904 181582 2916
rect 179564 2876 181582 2904
rect 179564 2864 179570 2876
rect 181576 2864 181582 2876
rect 181634 2864 181640 2916
rect 181714 2864 181720 2916
rect 181772 2904 181778 2916
rect 182680 2904 182686 2916
rect 181772 2876 182686 2904
rect 181772 2864 181778 2876
rect 182680 2864 182686 2876
rect 182738 2864 182744 2916
rect 187694 2864 187700 2916
rect 187752 2904 187758 2916
rect 189304 2904 189310 2916
rect 187752 2876 189310 2904
rect 187752 2864 187758 2876
rect 189304 2864 189310 2876
rect 189362 2864 189368 2916
rect 205634 2864 205640 2916
rect 205692 2904 205698 2916
rect 208072 2904 208078 2916
rect 205692 2876 208078 2904
rect 205692 2864 205698 2876
rect 208072 2864 208078 2876
rect 208130 2864 208136 2916
rect 211614 2864 211620 2916
rect 211672 2904 211678 2916
rect 213592 2904 213598 2916
rect 211672 2876 213598 2904
rect 211672 2864 211678 2876
rect 213592 2864 213598 2876
rect 213650 2864 213656 2916
rect 213730 2864 213736 2916
rect 213788 2904 213794 2916
rect 214696 2904 214702 2916
rect 213788 2876 214702 2904
rect 213788 2864 213794 2876
rect 214696 2864 214702 2876
rect 214754 2864 214760 2916
rect 214834 2864 214840 2916
rect 214892 2904 214898 2916
rect 215800 2904 215806 2916
rect 214892 2876 215806 2904
rect 214892 2864 214898 2876
rect 215800 2864 215806 2876
rect 215858 2864 215864 2916
rect 216674 2864 216680 2916
rect 216732 2904 216738 2916
rect 219112 2904 219118 2916
rect 216732 2876 219118 2904
rect 216732 2864 216738 2876
rect 219112 2864 219118 2876
rect 219170 2864 219176 2916
rect 220354 2864 220360 2916
rect 220412 2904 220418 2916
rect 221320 2904 221326 2916
rect 220412 2876 221326 2904
rect 220412 2864 220418 2876
rect 221320 2864 221326 2876
rect 221378 2864 221384 2916
rect 221458 2864 221464 2916
rect 221516 2904 221522 2916
rect 222424 2904 222430 2916
rect 221516 2876 222430 2904
rect 221516 2864 221522 2876
rect 222424 2864 222430 2876
rect 222482 2864 222488 2916
rect 222562 2864 222568 2916
rect 222620 2904 222626 2916
rect 224632 2904 224638 2916
rect 222620 2876 224638 2904
rect 222620 2864 222626 2876
rect 224632 2864 224638 2876
rect 224690 2864 224696 2916
rect 224770 2864 224776 2916
rect 224828 2904 224834 2916
rect 225736 2904 225742 2916
rect 224828 2876 225742 2904
rect 224828 2864 224834 2876
rect 225736 2864 225742 2876
rect 225794 2864 225800 2916
rect 226518 2864 226524 2916
rect 226576 2904 226582 2916
rect 227944 2904 227950 2916
rect 226576 2876 227950 2904
rect 226576 2864 226582 2876
rect 227944 2864 227950 2876
rect 228002 2864 228008 2916
rect 230566 2864 230572 2916
rect 230624 2904 230630 2916
rect 232360 2904 232366 2916
rect 230624 2876 232366 2904
rect 230624 2864 230630 2876
rect 232360 2864 232366 2876
rect 232418 2864 232424 2916
rect 232498 2864 232504 2916
rect 232556 2904 232562 2916
rect 233464 2904 233470 2916
rect 232556 2876 233470 2904
rect 232556 2864 232562 2876
rect 233464 2864 233470 2876
rect 233522 2864 233528 2916
rect 234706 2864 234712 2916
rect 234764 2904 234770 2916
rect 236776 2904 236782 2916
rect 234764 2876 236782 2904
rect 234764 2864 234770 2876
rect 236776 2864 236782 2876
rect 236834 2864 236840 2916
rect 242894 2864 242900 2916
rect 242952 2904 242958 2916
rect 246712 2904 246718 2916
rect 242952 2876 246718 2904
rect 242952 2864 242958 2876
rect 246712 2864 246718 2876
rect 246770 2864 246776 2916
rect 247586 2864 247592 2916
rect 247644 2904 247650 2916
rect 251128 2904 251134 2916
rect 247644 2876 251134 2904
rect 247644 2864 247650 2876
rect 251128 2864 251134 2876
rect 251186 2864 251192 2916
rect 253474 2864 253480 2916
rect 253532 2904 253538 2916
rect 256648 2904 256654 2916
rect 253532 2876 256654 2904
rect 253532 2864 253538 2876
rect 256648 2864 256654 2876
rect 256706 2864 256712 2916
rect 257062 2864 257068 2916
rect 257120 2904 257126 2916
rect 259960 2904 259966 2916
rect 257120 2876 259966 2904
rect 257120 2864 257126 2876
rect 259960 2864 259966 2876
rect 260018 2864 260024 2916
rect 261754 2864 261760 2916
rect 261812 2904 261818 2916
rect 264376 2904 264382 2916
rect 261812 2876 264382 2904
rect 261812 2864 261818 2876
rect 264376 2864 264382 2876
rect 264434 2864 264440 2916
rect 265342 2864 265348 2916
rect 265400 2904 265406 2916
rect 267688 2904 267694 2916
rect 265400 2876 267694 2904
rect 265400 2864 265406 2876
rect 267688 2864 267694 2876
rect 267746 2864 267752 2916
rect 267826 2864 267832 2916
rect 267884 2904 267890 2916
rect 269896 2904 269902 2916
rect 267884 2876 269902 2904
rect 267884 2864 267890 2876
rect 269896 2864 269902 2876
rect 269954 2864 269960 2916
rect 271230 2864 271236 2916
rect 271288 2904 271294 2916
rect 273208 2904 273214 2916
rect 271288 2876 273214 2904
rect 271288 2864 271294 2876
rect 273208 2864 273214 2876
rect 273266 2864 273272 2916
rect 273622 2864 273628 2916
rect 273680 2904 273686 2916
rect 275416 2904 275422 2916
rect 273680 2876 275422 2904
rect 273680 2864 273686 2876
rect 275416 2864 275422 2876
rect 275474 2864 275480 2916
rect 276014 2864 276020 2916
rect 276072 2904 276078 2916
rect 277624 2904 277630 2916
rect 276072 2876 277630 2904
rect 276072 2864 276078 2876
rect 277624 2864 277630 2876
rect 277682 2864 277688 2916
rect 278314 2864 278320 2916
rect 278372 2904 278378 2916
rect 279832 2904 279838 2916
rect 278372 2876 279838 2904
rect 278372 2864 278378 2876
rect 279832 2864 279838 2876
rect 279890 2864 279896 2916
rect 280706 2864 280712 2916
rect 280764 2904 280770 2916
rect 282040 2904 282046 2916
rect 280764 2876 282046 2904
rect 280764 2864 280770 2876
rect 282040 2864 282046 2876
rect 282098 2864 282104 2916
rect 283144 2864 283150 2916
rect 283202 2864 283208 2916
rect 286594 2864 286600 2916
rect 286652 2904 286658 2916
rect 287560 2904 287566 2916
rect 286652 2876 287566 2904
rect 286652 2864 286658 2876
rect 287560 2864 287566 2876
rect 287618 2864 287624 2916
rect 287790 2864 287796 2916
rect 287848 2904 287854 2916
rect 288664 2904 288670 2916
rect 287848 2876 288670 2904
rect 287848 2864 287854 2876
rect 288664 2864 288670 2876
rect 288722 2864 288728 2916
rect 293678 2864 293684 2916
rect 293736 2904 293742 2916
rect 294184 2904 294190 2916
rect 293736 2876 294190 2904
rect 293736 2864 293742 2876
rect 294184 2864 294190 2876
rect 294242 2864 294248 2916
rect 320680 2864 320686 2916
rect 320738 2904 320744 2916
rect 322106 2904 322112 2916
rect 320738 2876 322112 2904
rect 320738 2864 320744 2876
rect 322106 2864 322112 2876
rect 322164 2864 322170 2916
rect 322888 2864 322894 2916
rect 322946 2904 322952 2916
rect 324406 2904 324412 2916
rect 322946 2876 324412 2904
rect 322946 2864 322952 2876
rect 324406 2864 324412 2876
rect 324464 2864 324470 2916
rect 325096 2864 325102 2916
rect 325154 2904 325160 2916
rect 326798 2904 326804 2916
rect 325154 2876 326804 2904
rect 325154 2864 325160 2876
rect 326798 2864 326804 2876
rect 326856 2864 326862 2916
rect 329512 2864 329518 2916
rect 329570 2904 329576 2916
rect 331582 2904 331588 2916
rect 329570 2876 331588 2904
rect 329570 2864 329576 2876
rect 331582 2864 331588 2876
rect 331640 2864 331646 2916
rect 331720 2864 331726 2916
rect 331778 2904 331784 2916
rect 333790 2904 333796 2916
rect 331778 2876 333796 2904
rect 331778 2864 331784 2876
rect 333790 2864 333796 2876
rect 333848 2864 333854 2916
rect 335032 2864 335038 2916
rect 335090 2904 335096 2916
rect 336458 2904 336464 2916
rect 335090 2876 336464 2904
rect 335090 2864 335096 2876
rect 336458 2864 336464 2876
rect 336516 2864 336522 2916
rect 340552 2864 340558 2916
rect 340610 2904 340616 2916
rect 343358 2904 343364 2916
rect 340610 2876 343364 2904
rect 340610 2864 340616 2876
rect 343358 2864 343364 2876
rect 343416 2864 343422 2916
rect 346072 2864 346078 2916
rect 346130 2904 346136 2916
rect 347590 2904 347596 2916
rect 346130 2876 347596 2904
rect 346130 2864 346136 2876
rect 347590 2864 347596 2876
rect 347648 2864 347654 2916
rect 348280 2864 348286 2916
rect 348338 2904 348344 2916
rect 349890 2904 349896 2916
rect 348338 2876 349896 2904
rect 348338 2864 348344 2876
rect 349890 2864 349896 2876
rect 349948 2864 349954 2916
rect 352696 2864 352702 2916
rect 352754 2904 352760 2916
rect 355778 2904 355784 2916
rect 352754 2876 355784 2904
rect 352754 2864 352760 2876
rect 355778 2864 355784 2876
rect 355836 2864 355842 2916
rect 358216 2864 358222 2916
rect 358274 2904 358280 2916
rect 360102 2904 360108 2916
rect 358274 2876 360108 2904
rect 358274 2864 358280 2876
rect 360102 2864 360108 2876
rect 360160 2864 360166 2916
rect 362632 2864 362638 2916
rect 362690 2904 362696 2916
rect 363506 2904 363512 2916
rect 362690 2876 363512 2904
rect 362690 2864 362696 2876
rect 363506 2864 363512 2876
rect 363564 2864 363570 2916
rect 363736 2864 363742 2916
rect 363794 2904 363800 2916
rect 366174 2904 366180 2916
rect 363794 2876 366180 2904
rect 363794 2864 363800 2876
rect 366174 2864 366180 2876
rect 366232 2864 366238 2916
rect 369256 2864 369262 2916
rect 369314 2904 369320 2916
rect 370222 2904 370228 2916
rect 369314 2876 370228 2904
rect 369314 2864 369320 2876
rect 370222 2864 370228 2876
rect 370280 2864 370286 2916
rect 370360 2864 370366 2916
rect 370418 2904 370424 2916
rect 372706 2904 372712 2916
rect 370418 2876 372712 2904
rect 370418 2864 370424 2876
rect 372706 2864 372712 2876
rect 372764 2864 372770 2916
rect 373672 2864 373678 2916
rect 373730 2904 373736 2916
rect 375098 2904 375104 2916
rect 373730 2876 375104 2904
rect 373730 2864 373736 2876
rect 375098 2864 375104 2876
rect 375156 2864 375162 2916
rect 375880 2864 375886 2916
rect 375938 2904 375944 2916
rect 378502 2904 378508 2916
rect 375938 2876 378508 2904
rect 375938 2864 375944 2876
rect 378502 2864 378508 2876
rect 378560 2864 378566 2916
rect 379192 2864 379198 2916
rect 379250 2904 379256 2916
rect 380158 2904 380164 2916
rect 379250 2876 380164 2904
rect 379250 2864 379256 2876
rect 380158 2864 380164 2876
rect 380216 2864 380222 2916
rect 380296 2864 380302 2916
rect 380354 2904 380360 2916
rect 382274 2904 382280 2916
rect 380354 2876 382280 2904
rect 380354 2864 380360 2876
rect 382274 2864 382280 2876
rect 382332 2864 382338 2916
rect 386920 2864 386926 2916
rect 386978 2904 386984 2916
rect 387886 2904 387892 2916
rect 386978 2876 387892 2904
rect 386978 2864 386984 2876
rect 387886 2864 387892 2876
rect 387944 2864 387950 2916
rect 388024 2864 388030 2916
rect 388082 2904 388088 2916
rect 390646 2904 390652 2916
rect 388082 2876 390652 2904
rect 388082 2864 388088 2876
rect 390646 2864 390652 2876
rect 390704 2864 390710 2916
rect 391336 2864 391342 2916
rect 391394 2904 391400 2916
rect 394418 2904 394424 2916
rect 391394 2876 394424 2904
rect 391394 2864 391400 2876
rect 394418 2864 394424 2876
rect 394476 2864 394482 2916
rect 396856 2864 396862 2916
rect 396914 2904 396920 2916
rect 398742 2904 398748 2916
rect 396914 2876 398748 2904
rect 396914 2864 396920 2876
rect 398742 2864 398748 2876
rect 398800 2864 398806 2916
rect 399064 2864 399070 2916
rect 399122 2904 399128 2916
rect 401594 2904 401600 2916
rect 399122 2876 401600 2904
rect 399122 2864 399128 2876
rect 401594 2864 401600 2876
rect 401652 2864 401658 2916
rect 402376 2864 402382 2916
rect 402434 2904 402440 2916
rect 404262 2904 404268 2916
rect 402434 2876 404268 2904
rect 402434 2864 402440 2876
rect 404262 2864 404268 2876
rect 404320 2864 404326 2916
rect 406792 2864 406798 2916
rect 406850 2904 406856 2916
rect 407758 2904 407764 2916
rect 406850 2876 407764 2904
rect 406850 2864 406856 2876
rect 407758 2864 407764 2876
rect 407816 2864 407822 2916
rect 407896 2864 407902 2916
rect 407954 2904 407960 2916
rect 409782 2904 409788 2916
rect 407954 2876 409788 2904
rect 407954 2864 407960 2876
rect 409782 2864 409788 2876
rect 409840 2864 409846 2916
rect 415624 2864 415630 2916
rect 415682 2904 415688 2916
rect 423766 2904 423772 2916
rect 415682 2876 423772 2904
rect 415682 2864 415688 2876
rect 423766 2864 423772 2876
rect 423824 2864 423830 2916
rect 424456 2864 424462 2916
rect 424514 2904 424520 2916
rect 425422 2904 425428 2916
rect 424514 2876 425428 2904
rect 424514 2864 424520 2876
rect 425422 2864 425428 2876
rect 425480 2864 425486 2916
rect 425560 2864 425566 2916
rect 425618 2904 425624 2916
rect 428734 2904 428740 2916
rect 425618 2876 428740 2904
rect 425618 2864 425624 2876
rect 428734 2864 428740 2876
rect 428792 2864 428798 2916
rect 428872 2864 428878 2916
rect 428930 2904 428936 2916
rect 429838 2904 429844 2916
rect 428930 2876 429844 2904
rect 428930 2864 428936 2876
rect 429838 2864 429844 2876
rect 429896 2864 429902 2916
rect 429976 2864 429982 2916
rect 430034 2904 430040 2916
rect 433150 2904 433156 2916
rect 430034 2876 433156 2904
rect 430034 2864 430040 2876
rect 433150 2864 433156 2876
rect 433208 2864 433214 2916
rect 439912 2864 439918 2916
rect 439970 2904 439976 2916
rect 442902 2904 442908 2916
rect 439970 2876 442908 2904
rect 439970 2864 439976 2876
rect 442902 2864 442908 2876
rect 442960 2864 442966 2916
rect 450952 2864 450958 2916
rect 451010 2904 451016 2916
rect 452562 2904 452568 2916
rect 451010 2876 452568 2904
rect 451010 2864 451016 2876
rect 452562 2864 452568 2876
rect 452620 2864 452626 2916
rect 461992 2864 461998 2916
rect 462050 2904 462056 2916
rect 462050 2876 463004 2904
rect 462050 2864 462056 2876
rect 63494 2796 63500 2848
rect 63552 2836 63558 2848
rect 67864 2836 67870 2848
rect 63552 2808 67870 2836
rect 63552 2796 63558 2808
rect 67864 2796 67870 2808
rect 67922 2796 67928 2848
rect 73154 2796 73160 2848
rect 73212 2836 73218 2848
rect 75592 2836 75598 2848
rect 73212 2808 75598 2836
rect 73212 2796 73218 2808
rect 75592 2796 75598 2808
rect 75650 2796 75656 2848
rect 76834 2796 76840 2848
rect 76892 2836 76898 2848
rect 81112 2836 81118 2848
rect 76892 2808 81118 2836
rect 76892 2796 76898 2808
rect 81112 2796 81118 2808
rect 81170 2796 81176 2848
rect 100754 2796 100760 2848
rect 100812 2836 100818 2848
rect 103192 2836 103198 2848
rect 100812 2808 103198 2836
rect 100812 2796 100818 2808
rect 103192 2796 103198 2808
rect 103250 2796 103256 2848
rect 150434 2796 150440 2848
rect 150492 2836 150498 2848
rect 152872 2836 152878 2848
rect 150492 2808 152878 2836
rect 150492 2796 150498 2808
rect 152872 2796 152878 2808
rect 152930 2796 152936 2848
rect 204254 2796 204260 2848
rect 204312 2836 204318 2848
rect 206968 2836 206974 2848
rect 204312 2808 206974 2836
rect 204312 2796 204318 2808
rect 206968 2796 206974 2808
rect 207026 2796 207032 2848
rect 215294 2796 215300 2848
rect 215352 2836 215358 2848
rect 217962 2836 217968 2848
rect 215352 2808 217968 2836
rect 215352 2796 215358 2808
rect 217962 2796 217968 2808
rect 218020 2796 218026 2848
rect 218054 2796 218060 2848
rect 218112 2836 218118 2848
rect 220216 2836 220222 2848
rect 218112 2808 220222 2836
rect 218112 2796 218118 2808
rect 220216 2796 220222 2808
rect 220274 2796 220280 2848
rect 224954 2796 224960 2848
rect 225012 2836 225018 2848
rect 226840 2836 226846 2848
rect 225012 2808 226846 2836
rect 225012 2796 225018 2808
rect 226840 2796 226846 2808
rect 226898 2796 226904 2848
rect 249886 2796 249892 2848
rect 249944 2836 249950 2848
rect 253336 2836 253342 2848
rect 249944 2808 253342 2836
rect 249944 2796 249950 2808
rect 253336 2796 253342 2808
rect 253394 2796 253400 2848
rect 259454 2796 259460 2848
rect 259512 2836 259518 2848
rect 262168 2836 262174 2848
rect 259512 2808 262174 2836
rect 259512 2796 259518 2808
rect 262168 2796 262174 2808
rect 262226 2796 262232 2848
rect 266538 2796 266544 2848
rect 266596 2836 266602 2848
rect 268792 2836 268798 2848
rect 266596 2808 268798 2836
rect 266596 2796 266602 2808
rect 268792 2796 268798 2808
rect 268850 2796 268856 2848
rect 272426 2796 272432 2848
rect 272484 2836 272490 2848
rect 274312 2836 274318 2848
rect 272484 2808 274318 2836
rect 272484 2796 272490 2808
rect 274312 2796 274318 2808
rect 274370 2796 274376 2848
rect 274818 2796 274824 2848
rect 274876 2836 274882 2848
rect 276520 2836 276526 2848
rect 274876 2808 276526 2836
rect 274876 2796 274882 2808
rect 276520 2796 276526 2808
rect 276578 2796 276584 2848
rect 279510 2796 279516 2848
rect 279568 2836 279574 2848
rect 280936 2836 280942 2848
rect 279568 2808 280942 2836
rect 279568 2796 279574 2808
rect 280936 2796 280942 2808
rect 280994 2796 281000 2848
rect 281902 2796 281908 2848
rect 281960 2836 281966 2848
rect 283162 2836 283190 2864
rect 281960 2808 283190 2836
rect 281960 2796 281966 2808
rect 285398 2796 285404 2848
rect 285456 2836 285462 2848
rect 286456 2836 286462 2848
rect 285456 2808 286462 2836
rect 285456 2796 285462 2808
rect 286456 2796 286462 2808
rect 286514 2796 286520 2848
rect 316264 2796 316270 2848
rect 316322 2836 316328 2848
rect 317322 2836 317328 2848
rect 316322 2808 317328 2836
rect 316322 2796 316328 2808
rect 317322 2796 317328 2808
rect 317380 2796 317386 2848
rect 336136 2796 336142 2848
rect 336194 2836 336200 2848
rect 338666 2836 338672 2848
rect 336194 2808 338672 2836
rect 336194 2796 336200 2808
rect 338666 2796 338672 2808
rect 338724 2796 338730 2848
rect 342760 2796 342766 2848
rect 342818 2836 342824 2848
rect 345750 2836 345756 2848
rect 342818 2808 345756 2836
rect 342818 2796 342824 2808
rect 345750 2796 345756 2808
rect 345808 2796 345814 2848
rect 347176 2796 347182 2848
rect 347234 2836 347240 2848
rect 348786 2836 348792 2848
rect 347234 2808 348792 2836
rect 347234 2796 347240 2808
rect 348786 2796 348792 2808
rect 348844 2796 348850 2848
rect 349384 2796 349390 2848
rect 349442 2836 349448 2848
rect 352834 2836 352840 2848
rect 349442 2808 352840 2836
rect 349442 2796 349448 2808
rect 352834 2796 352840 2808
rect 352892 2796 352898 2848
rect 354904 2796 354910 2848
rect 354962 2836 354968 2848
rect 358722 2836 358728 2848
rect 354962 2808 358728 2836
rect 354962 2796 354968 2808
rect 358722 2796 358728 2808
rect 358780 2796 358786 2848
rect 359320 2796 359326 2848
rect 359378 2836 359384 2848
rect 362494 2836 362500 2848
rect 359378 2808 362500 2836
rect 359378 2796 359384 2808
rect 362494 2796 362500 2808
rect 362552 2796 362558 2848
rect 365944 2796 365950 2848
rect 366002 2836 366008 2848
rect 369762 2836 369768 2848
rect 366002 2808 369768 2836
rect 366002 2796 366008 2808
rect 369762 2796 369768 2808
rect 369820 2796 369826 2848
rect 374776 2796 374782 2848
rect 374834 2836 374840 2848
rect 376662 2836 376668 2848
rect 374834 2808 376668 2836
rect 374834 2796 374840 2808
rect 376662 2796 376668 2808
rect 376720 2796 376726 2848
rect 382504 2796 382510 2848
rect 382562 2836 382568 2848
rect 387702 2836 387708 2848
rect 382562 2808 387708 2836
rect 382562 2796 382568 2808
rect 387702 2796 387708 2808
rect 387760 2796 387766 2848
rect 393544 2796 393550 2848
rect 393602 2836 393608 2848
rect 396718 2836 396724 2848
rect 393602 2808 396724 2836
rect 393602 2796 393608 2808
rect 396718 2796 396724 2808
rect 396776 2796 396782 2848
rect 397960 2796 397966 2848
rect 398018 2836 398024 2848
rect 399846 2836 399852 2848
rect 398018 2808 399852 2836
rect 398018 2796 398024 2808
rect 399846 2796 399852 2808
rect 399904 2796 399910 2848
rect 403480 2796 403486 2848
rect 403538 2836 403544 2848
rect 407022 2836 407028 2848
rect 403538 2808 407028 2836
rect 403538 2796 403544 2808
rect 407022 2796 407028 2808
rect 407080 2796 407086 2848
rect 409000 2796 409006 2848
rect 409058 2836 409064 2848
rect 416590 2836 416596 2848
rect 409058 2808 416596 2836
rect 409058 2796 409064 2808
rect 416590 2796 416596 2808
rect 416648 2796 416654 2848
rect 432184 2796 432190 2848
rect 432242 2836 432248 2848
rect 438946 2836 438952 2848
rect 432242 2808 438952 2836
rect 432242 2796 432248 2808
rect 438946 2796 438952 2808
rect 439004 2796 439010 2848
rect 442120 2796 442126 2848
rect 442178 2836 442184 2848
rect 451182 2836 451188 2848
rect 442178 2808 451188 2836
rect 442178 2796 442184 2808
rect 451182 2796 451188 2808
rect 451240 2796 451246 2848
rect 452056 2796 452062 2848
rect 452114 2836 452120 2848
rect 462222 2836 462228 2848
rect 452114 2808 462228 2836
rect 452114 2796 452120 2808
rect 462222 2796 462228 2808
rect 462280 2796 462286 2848
rect 462976 2836 463004 2876
rect 463096 2864 463102 2916
rect 463154 2904 463160 2916
rect 464062 2904 464068 2916
rect 463154 2876 464068 2904
rect 463154 2864 463160 2876
rect 464062 2864 464068 2876
rect 464120 2864 464126 2916
rect 464200 2864 464206 2916
rect 464258 2904 464264 2916
rect 466178 2904 466184 2916
rect 464258 2876 466184 2904
rect 464258 2864 464264 2876
rect 466178 2864 466184 2876
rect 466236 2864 466242 2916
rect 476344 2864 476350 2916
rect 476402 2904 476408 2916
rect 478322 2904 478328 2916
rect 476402 2876 478328 2904
rect 476402 2864 476408 2876
rect 478322 2864 478328 2876
rect 478380 2864 478386 2916
rect 490696 2864 490702 2916
rect 490754 2904 490760 2916
rect 492582 2904 492588 2916
rect 490754 2876 492588 2904
rect 490754 2864 490760 2876
rect 492582 2864 492588 2876
rect 492640 2864 492646 2916
rect 506152 2864 506158 2916
rect 506210 2904 506216 2916
rect 507854 2904 507860 2916
rect 506210 2876 507860 2904
rect 506210 2864 506216 2876
rect 507854 2864 507860 2876
rect 507912 2864 507918 2916
rect 508360 2864 508366 2916
rect 508418 2904 508424 2916
rect 509970 2904 509976 2916
rect 508418 2876 509976 2904
rect 508418 2864 508424 2876
rect 509970 2864 509976 2876
rect 510028 2864 510034 2916
rect 523816 2864 523822 2916
rect 523874 2904 523880 2916
rect 525702 2904 525708 2916
rect 523874 2876 525708 2904
rect 523874 2864 523880 2876
rect 525702 2864 525708 2876
rect 525760 2864 525766 2916
rect 540376 2864 540382 2916
rect 540434 2904 540440 2916
rect 541342 2904 541348 2916
rect 540434 2876 541348 2904
rect 540434 2864 540440 2876
rect 541342 2864 541348 2876
rect 541400 2864 541406 2916
rect 541480 2864 541486 2916
rect 541538 2904 541544 2916
rect 556430 2904 556436 2916
rect 541538 2876 556436 2904
rect 541538 2864 541544 2876
rect 556430 2864 556436 2876
rect 556488 2864 556494 2916
rect 463602 2836 463608 2848
rect 462976 2808 463608 2836
rect 463602 2796 463608 2808
rect 463660 2796 463666 2848
rect 465304 2796 465310 2848
rect 465362 2836 465368 2848
rect 476942 2836 476948 2848
rect 465362 2808 476948 2836
rect 465362 2796 465368 2808
rect 476942 2796 476948 2808
rect 477000 2796 477006 2848
rect 478552 2796 478558 2848
rect 478610 2836 478616 2848
rect 488626 2836 488632 2848
rect 478610 2808 488632 2836
rect 478610 2796 478616 2808
rect 488626 2796 488632 2808
rect 488684 2796 488690 2848
rect 491800 2796 491806 2848
rect 491858 2836 491864 2848
rect 505370 2836 505376 2848
rect 491858 2808 505376 2836
rect 491858 2796 491864 2808
rect 505370 2796 505376 2808
rect 505428 2796 505434 2848
rect 509464 2796 509470 2848
rect 509522 2836 509528 2848
rect 524230 2836 524236 2848
rect 509522 2808 524236 2836
rect 509522 2796 509528 2808
rect 524230 2796 524236 2808
rect 524288 2796 524294 2848
rect 524920 2796 524926 2848
rect 524978 2836 524984 2848
rect 540790 2836 540796 2848
rect 524978 2808 540796 2836
rect 524978 2796 524984 2808
rect 540790 2796 540796 2808
rect 540848 2796 540854 2848
rect 28902 1300 28908 1352
rect 28960 1340 28966 1352
rect 28960 1312 31156 1340
rect 28960 1300 28966 1312
rect 23014 1232 23020 1284
rect 23072 1272 23078 1284
rect 23072 1244 31064 1272
rect 23072 1232 23078 1244
rect 17034 1096 17040 1148
rect 17092 1136 17098 1148
rect 17092 1108 26004 1136
rect 17092 1096 17098 1108
rect 18230 1028 18236 1080
rect 18288 1068 18294 1080
rect 25976 1068 26004 1108
rect 31036 1068 31064 1244
rect 31128 1136 31156 1312
rect 35986 1232 35992 1284
rect 36044 1272 36050 1284
rect 53466 1272 53472 1284
rect 36044 1244 53472 1272
rect 36044 1232 36050 1244
rect 53466 1232 53472 1244
rect 53524 1232 53530 1284
rect 31478 1164 31484 1216
rect 31536 1204 31542 1216
rect 44634 1204 44640 1216
rect 31536 1176 44640 1204
rect 31536 1164 31542 1176
rect 44634 1164 44640 1176
rect 44692 1164 44698 1216
rect 51350 1164 51356 1216
rect 51408 1204 51414 1216
rect 51408 1176 55214 1204
rect 51408 1164 51414 1176
rect 46842 1136 46848 1148
rect 31128 1108 46848 1136
rect 46842 1096 46848 1108
rect 46900 1096 46906 1148
rect 46952 1108 54800 1136
rect 41322 1068 41328 1080
rect 18288 1040 22692 1068
rect 25976 1040 26234 1068
rect 31036 1040 41328 1068
rect 18288 1028 18294 1040
rect 18874 960 18880 1012
rect 18932 1000 18938 1012
rect 22554 1000 22560 1012
rect 18932 972 22560 1000
rect 18932 960 18938 972
rect 22554 960 22560 972
rect 22612 960 22618 1012
rect 22664 1000 22692 1040
rect 26206 1000 26234 1040
rect 41322 1028 41328 1040
rect 41380 1028 41386 1080
rect 46658 1028 46664 1080
rect 46716 1068 46722 1080
rect 46952 1068 46980 1108
rect 46716 1040 46980 1068
rect 46716 1028 46722 1040
rect 35802 1000 35808 1012
rect 22664 972 26004 1000
rect 26206 972 35808 1000
rect 21174 892 21180 944
rect 21232 932 21238 944
rect 25866 932 25872 944
rect 21232 904 25872 932
rect 21232 892 21238 904
rect 25866 892 25872 904
rect 25924 892 25930 944
rect 25976 932 26004 972
rect 35802 960 35808 972
rect 35860 960 35866 1012
rect 40678 960 40684 1012
rect 40736 1000 40742 1012
rect 40736 972 45554 1000
rect 40736 960 40742 972
rect 36906 932 36912 944
rect 25976 904 36912 932
rect 36906 892 36912 904
rect 36964 892 36970 944
rect 45526 932 45554 972
rect 47210 960 47216 1012
rect 47268 1000 47274 1012
rect 54570 1000 54576 1012
rect 47268 972 54576 1000
rect 47268 960 47274 972
rect 54570 960 54576 972
rect 54628 960 54634 1012
rect 54772 1000 54800 1108
rect 55186 1068 55214 1176
rect 65518 1164 65524 1216
rect 65576 1204 65582 1216
rect 118602 1204 118608 1216
rect 65576 1176 74534 1204
rect 65576 1164 65582 1176
rect 58434 1096 58440 1148
rect 58492 1136 58498 1148
rect 71774 1136 71780 1148
rect 58492 1108 71780 1136
rect 58492 1096 58498 1108
rect 71774 1096 71780 1108
rect 71832 1096 71838 1148
rect 74506 1136 74534 1176
rect 111444 1176 118608 1204
rect 76834 1136 76840 1148
rect 74506 1108 76840 1136
rect 76834 1096 76840 1108
rect 76892 1096 76898 1148
rect 77386 1096 77392 1148
rect 77444 1136 77450 1148
rect 88150 1136 88156 1148
rect 77444 1108 88156 1136
rect 77444 1096 77450 1108
rect 88150 1096 88156 1108
rect 88208 1096 88214 1148
rect 63494 1068 63500 1080
rect 55186 1040 63500 1068
rect 63494 1028 63500 1040
rect 63552 1028 63558 1080
rect 69106 1028 69112 1080
rect 69164 1068 69170 1080
rect 80146 1068 80152 1080
rect 69164 1040 80152 1068
rect 69164 1028 69170 1040
rect 80146 1028 80152 1040
rect 80204 1028 80210 1080
rect 97442 1028 97448 1080
rect 97500 1068 97506 1080
rect 110874 1068 110880 1080
rect 97500 1040 110880 1068
rect 97500 1028 97506 1040
rect 110874 1028 110880 1040
rect 110932 1028 110938 1080
rect 63402 1000 63408 1012
rect 54772 972 63408 1000
rect 63402 960 63408 972
rect 63460 960 63466 1012
rect 71498 960 71504 1012
rect 71556 1000 71562 1012
rect 85390 1000 85396 1012
rect 71556 972 85396 1000
rect 71556 960 71562 972
rect 85390 960 85396 972
rect 85448 960 85454 1012
rect 91554 960 91560 1012
rect 91612 1000 91618 1012
rect 102226 1000 102232 1012
rect 91612 972 102232 1000
rect 91612 960 91618 972
rect 102226 960 102232 972
rect 102284 960 102290 1012
rect 57882 932 57888 944
rect 45526 904 57888 932
rect 57882 892 57888 904
rect 57940 892 57946 944
rect 59630 892 59636 944
rect 59688 932 59694 944
rect 73154 932 73160 944
rect 59688 904 73160 932
rect 59688 892 59694 904
rect 73154 892 73160 904
rect 73212 892 73218 944
rect 83274 892 83280 944
rect 83332 932 83338 944
rect 83332 904 84194 932
rect 83332 892 83338 904
rect 11146 824 11152 876
rect 11204 864 11210 876
rect 30282 864 30288 876
rect 11204 836 30288 864
rect 11204 824 11210 836
rect 30282 824 30288 836
rect 30340 824 30346 876
rect 30374 824 30380 876
rect 30432 864 30438 876
rect 47946 864 47952 876
rect 30432 836 47952 864
rect 30432 824 30438 836
rect 47946 824 47952 836
rect 48004 824 48010 876
rect 59170 864 59176 876
rect 52472 836 59176 864
rect 12342 756 12348 808
rect 12400 796 12406 808
rect 31386 796 31392 808
rect 12400 768 31392 796
rect 12400 756 12406 768
rect 31386 756 31392 768
rect 31444 756 31450 808
rect 34790 756 34796 808
rect 34848 796 34854 808
rect 52362 796 52368 808
rect 34848 768 52368 796
rect 34848 756 34854 768
rect 52362 756 52368 768
rect 52420 756 52426 808
rect 13538 688 13544 740
rect 13596 728 13602 740
rect 32490 728 32496 740
rect 13596 700 32496 728
rect 13596 688 13602 700
rect 32490 688 32496 700
rect 32548 688 32554 740
rect 41874 688 41880 740
rect 41932 728 41938 740
rect 41932 700 45554 728
rect 41932 688 41938 700
rect 5258 620 5264 672
rect 5316 660 5322 672
rect 24762 660 24768 672
rect 5316 632 24768 660
rect 5316 620 5322 632
rect 24762 620 24768 632
rect 24820 620 24826 672
rect 42426 660 42432 672
rect 24872 632 42432 660
rect 6454 552 6460 604
rect 6512 592 6518 604
rect 21174 592 21180 604
rect 6512 564 21180 592
rect 6512 552 6518 564
rect 21174 552 21180 564
rect 21232 552 21238 604
rect 24210 552 24216 604
rect 24268 592 24274 604
rect 24872 592 24900 632
rect 42426 620 42432 632
rect 42484 620 42490 672
rect 43530 660 43536 672
rect 42536 632 43536 660
rect 24268 564 24900 592
rect 24268 552 24274 564
rect 25314 552 25320 604
rect 25372 592 25378 604
rect 42536 592 42564 632
rect 43530 620 43536 632
rect 43588 620 43594 672
rect 45526 660 45554 700
rect 47854 688 47860 740
rect 47912 728 47918 740
rect 52472 728 52500 836
rect 59170 824 59176 836
rect 59228 824 59234 876
rect 60826 824 60832 876
rect 60884 864 60890 876
rect 60884 836 69060 864
rect 60884 824 60890 836
rect 53742 756 53748 808
rect 53800 796 53806 808
rect 67634 796 67640 808
rect 53800 768 67640 796
rect 53800 756 53806 768
rect 67634 756 67640 768
rect 67692 756 67698 808
rect 47912 700 52500 728
rect 47912 688 47918 700
rect 52546 688 52552 740
rect 52604 728 52610 740
rect 68922 728 68928 740
rect 52604 700 68928 728
rect 52604 688 52610 700
rect 68922 688 68928 700
rect 68980 688 68986 740
rect 58986 660 58992 672
rect 45526 632 58992 660
rect 58986 620 58992 632
rect 59044 620 59050 672
rect 64322 620 64328 672
rect 64380 660 64386 672
rect 69032 660 69060 836
rect 76926 824 76932 876
rect 76984 864 76990 876
rect 82170 864 82176 876
rect 76984 836 82176 864
rect 76984 824 76990 836
rect 82170 824 82176 836
rect 82228 824 82234 876
rect 84166 864 84194 904
rect 86862 892 86868 944
rect 86920 932 86926 944
rect 97994 932 98000 944
rect 86920 904 98000 932
rect 86920 892 86926 904
rect 97994 892 98000 904
rect 98052 892 98058 944
rect 100754 932 100760 944
rect 98196 904 100760 932
rect 95694 864 95700 876
rect 84166 836 95700 864
rect 95694 824 95700 836
rect 95752 824 95758 876
rect 98196 864 98224 904
rect 100754 892 100760 904
rect 100812 892 100818 944
rect 105722 892 105728 944
rect 105780 932 105786 944
rect 111444 932 111472 1176
rect 118602 1164 118608 1176
rect 118660 1164 118666 1216
rect 537110 1164 537116 1216
rect 537168 1204 537174 1216
rect 553762 1204 553768 1216
rect 537168 1176 553768 1204
rect 537168 1164 537174 1176
rect 553762 1164 553768 1176
rect 553820 1164 553826 1216
rect 114738 1136 114744 1148
rect 105780 904 111472 932
rect 111536 1108 114744 1136
rect 105780 892 105786 904
rect 96080 836 98224 864
rect 72602 756 72608 808
rect 72660 796 72666 808
rect 86770 796 86776 808
rect 72660 768 86776 796
rect 72660 756 72666 768
rect 86770 756 86776 768
rect 86828 756 86834 808
rect 89162 756 89168 808
rect 89220 796 89226 808
rect 96080 796 96108 836
rect 99834 824 99840 876
rect 99892 864 99898 876
rect 110414 864 110420 876
rect 99892 836 110420 864
rect 99892 824 99898 836
rect 110414 824 110420 836
rect 110472 824 110478 876
rect 102042 796 102048 808
rect 89220 768 96108 796
rect 96172 768 102048 796
rect 89220 756 89226 768
rect 70302 688 70308 740
rect 70360 728 70366 740
rect 85482 728 85488 740
rect 70360 700 85488 728
rect 70360 688 70366 700
rect 85482 688 85488 700
rect 85540 688 85546 740
rect 87966 688 87972 740
rect 88024 728 88030 740
rect 96172 728 96200 768
rect 102042 756 102048 768
rect 102100 756 102106 808
rect 105998 756 106004 808
rect 106056 796 106062 808
rect 107746 796 107752 808
rect 106056 768 107752 796
rect 106056 756 106062 768
rect 107746 756 107752 768
rect 107804 756 107810 808
rect 88024 700 96200 728
rect 88024 688 88030 700
rect 96246 688 96252 740
rect 96304 728 96310 740
rect 96304 700 101260 728
rect 96304 688 96310 700
rect 75454 660 75460 672
rect 64380 632 67036 660
rect 69032 632 75460 660
rect 64380 620 64386 632
rect 25372 564 42564 592
rect 25372 552 25378 564
rect 43070 552 43076 604
rect 43128 592 43134 604
rect 60090 592 60096 604
rect 43128 564 60096 592
rect 43128 552 43134 564
rect 60090 552 60096 564
rect 60148 552 60154 604
rect 62022 552 62028 604
rect 62080 592 62086 604
rect 67008 592 67036 632
rect 75454 620 75460 632
rect 75512 620 75518 672
rect 76190 620 76196 672
rect 76248 660 76254 672
rect 91002 660 91008 672
rect 76248 632 91008 660
rect 76248 620 76254 632
rect 91002 620 91008 632
rect 91060 620 91066 672
rect 95142 620 95148 672
rect 95200 660 95206 672
rect 95200 632 101168 660
rect 95200 620 95206 632
rect 62080 564 66944 592
rect 67008 564 77892 592
rect 62080 552 62086 564
rect 14550 484 14556 536
rect 14608 524 14614 536
rect 33410 524 33416 536
rect 14608 496 33416 524
rect 14608 484 14614 496
rect 33410 484 33416 496
rect 33468 484 33474 536
rect 36998 484 37004 536
rect 37056 524 37062 536
rect 47210 524 47216 536
rect 37056 496 47216 524
rect 37056 484 37062 496
rect 47210 484 47216 496
rect 47268 484 47274 536
rect 49142 524 49148 536
rect 47320 496 49148 524
rect 7834 416 7840 468
rect 7892 456 7898 468
rect 26970 456 26976 468
rect 7892 428 26976 456
rect 7892 416 7898 428
rect 26970 416 26976 428
rect 27028 416 27034 468
rect 31110 416 31116 468
rect 31168 456 31174 468
rect 47320 456 47348 496
rect 49142 484 49148 496
rect 49200 484 49206 536
rect 66916 524 66944 564
rect 77754 524 77760 536
rect 66916 496 77760 524
rect 77754 484 77760 496
rect 77812 484 77818 536
rect 31168 428 47348 456
rect 31168 416 31174 428
rect 48774 416 48780 468
rect 48832 456 48838 468
rect 65702 456 65708 468
rect 48832 428 65708 456
rect 48832 416 48838 428
rect 65702 416 65708 428
rect 65760 416 65766 468
rect 66898 416 66904 468
rect 66956 456 66962 468
rect 76926 456 76932 468
rect 66956 428 76932 456
rect 66956 416 66962 428
rect 76926 416 76932 428
rect 76984 416 76990 468
rect 77864 456 77892 564
rect 79686 552 79692 604
rect 79744 552 79750 604
rect 82078 552 82084 604
rect 82136 592 82142 604
rect 96522 592 96528 604
rect 82136 564 96528 592
rect 82136 552 82142 564
rect 96522 552 96528 564
rect 96580 552 96586 604
rect 101030 552 101036 604
rect 101088 552 101094 604
rect 79704 524 79732 552
rect 92474 524 92480 536
rect 79704 496 92480 524
rect 92474 484 92480 496
rect 92532 484 92538 536
rect 79962 456 79968 468
rect 77864 428 79968 456
rect 79962 416 79968 428
rect 80020 416 80026 468
rect 84654 416 84660 468
rect 84712 456 84718 468
rect 98822 456 98828 468
rect 84712 428 98828 456
rect 84712 416 84718 428
rect 98822 416 98828 428
rect 98880 416 98886 468
rect 101048 456 101076 552
rect 101140 524 101168 632
rect 101232 592 101260 700
rect 103330 688 103336 740
rect 103388 728 103394 740
rect 111536 728 111564 1108
rect 114738 1096 114744 1108
rect 114796 1096 114802 1148
rect 541342 1096 541348 1148
rect 541400 1136 541406 1148
rect 557350 1136 557356 1148
rect 541400 1108 557356 1136
rect 541400 1096 541406 1108
rect 557350 1096 557356 1108
rect 557408 1096 557414 1148
rect 111610 1028 111616 1080
rect 111668 1068 111674 1080
rect 111668 1040 118694 1068
rect 111668 1028 111674 1040
rect 117314 932 117320 944
rect 103388 700 111564 728
rect 112548 904 117320 932
rect 103388 688 103394 700
rect 101306 620 101312 672
rect 101364 660 101370 672
rect 107562 660 107568 672
rect 101364 632 107568 660
rect 101364 620 101370 632
rect 107562 620 107568 632
rect 107620 620 107626 672
rect 112548 660 112576 904
rect 117314 892 117320 904
rect 117372 892 117378 944
rect 118666 932 118694 1040
rect 509970 1028 509976 1080
rect 510028 1068 510034 1080
rect 523034 1068 523040 1080
rect 510028 1040 523040 1068
rect 510028 1028 510034 1040
rect 523034 1028 523040 1040
rect 523092 1028 523098 1080
rect 525702 1028 525708 1080
rect 525760 1068 525766 1080
rect 539594 1068 539600 1080
rect 525760 1040 539600 1068
rect 525760 1028 525766 1040
rect 539594 1028 539600 1040
rect 539652 1028 539658 1080
rect 548150 1028 548156 1080
rect 548208 1068 548214 1080
rect 565630 1068 565636 1080
rect 548208 1040 565636 1068
rect 548208 1028 548214 1040
rect 565630 1028 565636 1040
rect 565688 1028 565694 1080
rect 143442 960 143448 1012
rect 143500 1000 143506 1012
rect 149054 1000 149060 1012
rect 143500 972 149060 1000
rect 143500 960 143506 972
rect 149054 960 149060 972
rect 149112 960 149118 1012
rect 470870 960 470876 1012
rect 470928 1000 470934 1012
rect 482830 1000 482836 1012
rect 470928 972 482836 1000
rect 470928 960 470934 972
rect 482830 960 482836 972
rect 482888 960 482894 1012
rect 487430 960 487436 1012
rect 487488 1000 487494 1012
rect 500586 1000 500592 1012
rect 487488 972 500592 1000
rect 487488 960 487494 972
rect 500586 960 500592 972
rect 500644 960 500650 1012
rect 501782 960 501788 1012
rect 501840 1000 501846 1012
rect 506106 1000 506112 1012
rect 501840 972 506112 1000
rect 501840 960 501846 972
rect 506106 960 506112 972
rect 506164 960 506170 1012
rect 507854 960 507860 1012
rect 507912 1000 507918 1012
rect 507912 972 518894 1000
rect 507912 960 507918 972
rect 120074 932 120080 944
rect 118666 904 120080 932
rect 120074 892 120080 904
rect 120132 892 120138 944
rect 127526 892 127532 944
rect 127584 932 127590 944
rect 133230 932 133236 944
rect 127584 904 133236 932
rect 127584 892 127590 904
rect 133230 892 133236 904
rect 133288 892 133294 944
rect 135254 892 135260 944
rect 135312 932 135318 944
rect 144178 932 144184 944
rect 135312 904 144184 932
rect 135312 892 135318 904
rect 144178 892 144184 904
rect 144236 892 144242 944
rect 148318 892 148324 944
rect 148376 932 148382 944
rect 155954 932 155960 944
rect 148376 904 155960 932
rect 148376 892 148382 904
rect 155954 892 155960 904
rect 156012 892 156018 944
rect 190822 892 190828 944
rect 190880 932 190886 944
rect 198090 932 198096 944
rect 190880 904 198096 932
rect 190880 892 190886 904
rect 198090 892 198096 904
rect 198148 892 198154 944
rect 466178 892 466184 944
rect 466236 932 466242 944
rect 475746 932 475752 944
rect 466236 904 475752 932
rect 466236 892 466242 904
rect 475746 892 475752 904
rect 475804 892 475810 944
rect 478322 892 478328 944
rect 478380 932 478386 944
rect 488810 932 488816 944
rect 478380 904 488816 932
rect 478380 892 478386 904
rect 488810 892 488816 904
rect 488868 892 488874 944
rect 492582 892 492588 944
rect 492640 932 492646 944
rect 492640 904 503944 932
rect 492640 892 492646 904
rect 115198 824 115204 876
rect 115256 864 115262 876
rect 125134 864 125140 876
rect 115256 836 125140 864
rect 115256 824 115262 836
rect 125134 824 125140 836
rect 125192 824 125198 876
rect 128170 824 128176 876
rect 128228 864 128234 876
rect 136634 864 136640 876
rect 128228 836 136640 864
rect 128228 824 128234 836
rect 136634 824 136640 836
rect 136692 824 136698 876
rect 140038 824 140044 876
rect 140096 864 140102 876
rect 150618 864 150624 876
rect 140096 836 150624 864
rect 140096 824 140102 836
rect 150618 824 150624 836
rect 150676 824 150682 876
rect 161474 824 161480 876
rect 161532 864 161538 876
rect 169570 864 169576 876
rect 161532 836 169576 864
rect 161532 824 161538 836
rect 169570 824 169576 836
rect 169628 824 169634 876
rect 183738 824 183744 876
rect 183796 864 183802 876
rect 191466 864 191472 876
rect 183796 836 191472 864
rect 183796 824 183802 836
rect 191466 824 191472 836
rect 191524 824 191530 876
rect 210970 824 210976 876
rect 211028 864 211034 876
rect 216858 864 216864 876
rect 211028 836 216864 864
rect 211028 824 211034 836
rect 216858 824 216864 836
rect 216916 824 216922 876
rect 433058 824 433064 876
rect 433116 864 433122 876
rect 433242 864 433248 876
rect 433116 836 433248 864
rect 433116 824 433122 836
rect 433242 824 433248 836
rect 433300 824 433306 876
rect 464062 824 464068 876
rect 464120 864 464126 876
rect 474550 864 474556 876
rect 464120 836 474556 864
rect 464120 824 464126 836
rect 474550 824 474556 836
rect 474608 824 474614 876
rect 475286 824 475292 876
rect 475344 864 475350 876
rect 487614 864 487620 876
rect 475344 836 487620 864
rect 475344 824 475350 836
rect 487614 824 487620 836
rect 487672 824 487678 876
rect 492950 824 492956 876
rect 493008 864 493014 876
rect 503916 864 503944 904
rect 503990 892 503996 944
rect 504048 932 504054 944
rect 518250 932 518256 944
rect 504048 904 518256 932
rect 504048 892 504054 904
rect 518250 892 518256 904
rect 518308 892 518314 944
rect 518866 932 518894 972
rect 520550 960 520556 1012
rect 520608 1000 520614 1012
rect 536098 1000 536104 1012
rect 520608 972 536104 1000
rect 520608 960 520614 972
rect 536098 960 536104 972
rect 536156 960 536162 1012
rect 547046 960 547052 1012
rect 547104 1000 547110 1012
rect 564434 1000 564440 1012
rect 547104 972 564440 1000
rect 547104 960 547110 972
rect 564434 960 564440 972
rect 564492 960 564498 1012
rect 520734 932 520740 944
rect 518866 904 520740 932
rect 520734 892 520740 904
rect 520792 892 520798 944
rect 526070 892 526076 944
rect 526128 932 526134 944
rect 541986 932 541992 944
rect 526128 904 541992 932
rect 526128 892 526134 904
rect 541986 892 541992 904
rect 542044 892 542050 944
rect 545942 892 545948 944
rect 546000 932 546006 944
rect 563238 932 563244 944
rect 546000 904 563244 932
rect 546000 892 546006 904
rect 563238 892 563244 904
rect 563296 892 563302 944
rect 504174 864 504180 876
rect 493008 836 503760 864
rect 503916 836 504180 864
rect 493008 824 493014 836
rect 112806 756 112812 808
rect 112864 796 112870 808
rect 112864 768 116624 796
rect 112864 756 112870 768
rect 107672 632 112576 660
rect 113836 632 116532 660
rect 105998 592 106004 604
rect 101232 564 106004 592
rect 105998 552 106004 564
rect 106056 552 106062 604
rect 101140 496 106136 524
rect 101048 428 106044 456
rect 8938 348 8944 400
rect 8996 388 9002 400
rect 8996 360 21312 388
rect 8996 348 9002 360
rect 9766 280 9772 332
rect 9824 320 9830 332
rect 21174 320 21180 332
rect 9824 292 21180 320
rect 9824 280 9830 292
rect 21174 280 21180 292
rect 21232 280 21238 332
rect 1486 212 1492 264
rect 1544 252 1550 264
rect 21284 252 21312 360
rect 21358 348 21364 400
rect 21416 388 21422 400
rect 21416 360 21496 388
rect 21416 348 21422 360
rect 21468 320 21496 360
rect 26326 348 26332 400
rect 26384 388 26390 400
rect 31478 388 31484 400
rect 26384 360 31484 388
rect 26384 348 26390 360
rect 31478 348 31484 360
rect 31536 348 31542 400
rect 32214 348 32220 400
rect 32272 388 32278 400
rect 49970 388 49976 400
rect 32272 360 49976 388
rect 32272 348 32278 360
rect 49970 348 49976 360
rect 50028 348 50034 400
rect 55122 348 55128 400
rect 55180 388 55186 400
rect 71130 388 71136 400
rect 55180 360 71136 388
rect 55180 348 55186 360
rect 71130 348 71136 360
rect 71188 348 71194 400
rect 78398 348 78404 400
rect 78456 388 78462 400
rect 78456 360 88932 388
rect 78456 348 78462 360
rect 29178 320 29184 332
rect 21468 292 29184 320
rect 29178 280 29184 292
rect 29236 280 29242 332
rect 33778 280 33784 332
rect 33836 320 33842 332
rect 51166 320 51172 332
rect 33836 292 51172 320
rect 33836 280 33842 292
rect 51166 280 51172 292
rect 51224 280 51230 332
rect 56226 280 56232 332
rect 56284 320 56290 332
rect 72234 320 72240 332
rect 56284 292 72240 320
rect 56284 280 56290 292
rect 72234 280 72240 292
rect 72292 280 72298 332
rect 73614 280 73620 332
rect 73672 320 73678 332
rect 88794 320 88800 332
rect 73672 292 88800 320
rect 73672 280 73678 292
rect 88794 280 88800 292
rect 88852 280 88858 332
rect 88904 320 88932 360
rect 92566 348 92572 400
rect 92624 388 92630 400
rect 105538 388 105544 400
rect 92624 360 105544 388
rect 92624 348 92630 360
rect 105538 348 105544 360
rect 105596 348 105602 400
rect 93210 320 93216 332
rect 88904 292 93216 320
rect 93210 280 93216 292
rect 93268 280 93274 332
rect 94130 280 94136 332
rect 94188 320 94194 332
rect 101306 320 101312 332
rect 94188 292 101312 320
rect 94188 280 94194 292
rect 101306 280 101312 292
rect 101364 280 101370 332
rect 106016 320 106044 428
rect 106108 388 106136 496
rect 106734 484 106740 536
rect 106792 524 106798 536
rect 107672 524 107700 632
rect 108114 552 108120 604
rect 108172 592 108178 604
rect 113836 592 113864 632
rect 108172 564 113864 592
rect 108172 552 108178 564
rect 114186 524 114192 536
rect 106792 496 107700 524
rect 108960 496 114192 524
rect 106792 484 106798 496
rect 108666 388 108672 400
rect 106108 360 108672 388
rect 108666 348 108672 360
rect 108724 348 108730 400
rect 108960 320 108988 496
rect 114186 484 114192 496
rect 114244 484 114250 536
rect 116504 524 116532 632
rect 116596 592 116624 768
rect 123478 756 123484 808
rect 123536 796 123542 808
rect 123536 768 127756 796
rect 123536 756 123542 768
rect 117590 688 117596 740
rect 117648 728 117654 740
rect 127618 728 127624 740
rect 117648 700 127624 728
rect 117648 688 117654 700
rect 127618 688 127624 700
rect 127676 688 127682 740
rect 127728 728 127756 768
rect 129366 756 129372 808
rect 129424 796 129430 808
rect 140682 796 140688 808
rect 129424 768 140688 796
rect 129424 756 129430 768
rect 140682 756 140688 768
rect 140740 756 140746 808
rect 141234 756 141240 808
rect 141292 796 141298 808
rect 143442 796 143448 808
rect 141292 768 143448 796
rect 141292 756 141298 768
rect 143442 756 143448 768
rect 143500 756 143506 808
rect 143534 756 143540 808
rect 143592 796 143598 808
rect 153930 796 153936 808
rect 143592 768 153936 796
rect 143592 756 143598 768
rect 153930 756 153936 768
rect 153988 756 153994 808
rect 164878 756 164884 808
rect 164936 796 164942 808
rect 173802 796 173808 808
rect 164936 768 173808 796
rect 164936 756 164942 768
rect 173802 756 173808 768
rect 173860 756 173866 808
rect 184934 756 184940 808
rect 184992 796 184998 808
rect 192570 796 192576 808
rect 184992 768 192576 796
rect 184992 756 184998 768
rect 192570 756 192576 768
rect 192628 756 192634 808
rect 193214 756 193220 808
rect 193272 796 193278 808
rect 200298 796 200304 808
rect 193272 768 200304 796
rect 193272 756 193278 768
rect 200298 756 200304 768
rect 200356 756 200362 808
rect 203886 756 203892 808
rect 203944 796 203950 808
rect 210234 796 210240 808
rect 203944 768 210240 796
rect 203944 756 203950 768
rect 210234 756 210240 768
rect 210292 756 210298 808
rect 214466 756 214472 808
rect 214524 796 214530 808
rect 218054 796 218060 808
rect 214524 768 218060 796
rect 214524 756 214530 768
rect 218054 756 218060 768
rect 218112 756 218118 808
rect 223942 756 223948 808
rect 224000 796 224006 808
rect 229002 796 229008 808
rect 224000 768 229008 796
rect 224000 756 224006 768
rect 229002 756 229008 768
rect 229060 756 229066 808
rect 229830 756 229836 808
rect 229888 796 229894 808
rect 234522 796 234528 808
rect 229888 768 234528 796
rect 229888 756 229894 768
rect 234522 756 234528 768
rect 234580 756 234586 808
rect 351638 756 351644 808
rect 351696 796 351702 808
rect 355226 796 355232 808
rect 351696 768 355232 796
rect 351696 756 351702 768
rect 355226 756 355232 768
rect 355284 756 355290 808
rect 367002 756 367008 808
rect 367060 796 367066 808
rect 371694 796 371700 808
rect 367060 768 371700 796
rect 367060 756 367066 768
rect 371694 756 371700 768
rect 371752 756 371758 808
rect 378042 756 378048 808
rect 378100 796 378106 808
rect 383562 796 383568 808
rect 378100 768 383568 796
rect 378100 756 378106 768
rect 383562 756 383568 768
rect 383620 756 383626 808
rect 385862 756 385868 808
rect 385920 796 385926 808
rect 391842 796 391848 808
rect 385920 768 391848 796
rect 385920 756 385926 768
rect 391842 756 391848 768
rect 391900 756 391906 808
rect 394510 756 394516 808
rect 394568 796 394574 808
rect 401318 796 401324 808
rect 394568 768 401324 796
rect 394568 756 394574 768
rect 401318 756 401324 768
rect 401376 756 401382 808
rect 404630 756 404636 808
rect 404688 796 404694 808
rect 411898 796 411904 808
rect 404688 768 411904 796
rect 404688 756 404694 768
rect 411898 756 411904 768
rect 411956 756 411962 808
rect 416682 756 416688 808
rect 416740 796 416746 808
rect 424962 796 424968 808
rect 416740 768 424968 796
rect 416740 756 416746 768
rect 424962 756 424968 768
rect 425020 756 425026 808
rect 433150 756 433156 808
rect 433208 796 433214 808
rect 439130 796 439136 808
rect 433208 768 439136 796
rect 433208 756 433214 768
rect 439130 756 439136 768
rect 439188 756 439194 808
rect 443270 756 443276 808
rect 443328 796 443334 808
rect 451090 796 451096 808
rect 443328 768 451096 796
rect 443328 756 443334 768
rect 451090 756 451096 768
rect 451148 756 451154 808
rect 471054 796 471060 808
rect 462976 768 471060 796
rect 135162 728 135168 740
rect 127728 700 135168 728
rect 135162 688 135168 700
rect 135220 688 135226 740
rect 144730 688 144736 740
rect 144788 728 144794 740
rect 153378 728 153384 740
rect 144788 700 153384 728
rect 144788 688 144794 700
rect 153378 688 153384 700
rect 153436 688 153442 740
rect 166166 688 166172 740
rect 166224 728 166230 740
rect 172974 728 172980 740
rect 166224 700 172980 728
rect 166224 688 166230 700
rect 172974 688 172980 700
rect 173032 688 173038 740
rect 173158 688 173164 740
rect 173216 728 173222 740
rect 179506 728 179512 740
rect 173216 700 179512 728
rect 173216 688 173222 700
rect 179506 688 179512 700
rect 179564 688 179570 740
rect 181438 688 181444 740
rect 181496 728 181502 740
rect 187694 728 187700 740
rect 181496 700 187700 728
rect 181496 688 181502 700
rect 187694 688 187700 700
rect 187752 688 187758 740
rect 190362 728 190368 740
rect 187804 700 190368 728
rect 118786 620 118792 672
rect 118844 660 118850 672
rect 130746 660 130752 672
rect 118844 632 130752 660
rect 118844 620 118850 632
rect 130746 620 130752 632
rect 130804 620 130810 672
rect 136450 620 136456 672
rect 136508 660 136514 672
rect 147306 660 147312 672
rect 136508 632 147312 660
rect 136508 620 136514 632
rect 147306 620 147312 632
rect 147364 620 147370 672
rect 149514 620 149520 672
rect 149572 660 149578 672
rect 159450 660 159456 672
rect 149572 632 159456 660
rect 149572 620 149578 632
rect 159450 620 159456 632
rect 159508 620 159514 672
rect 160094 620 160100 672
rect 160152 660 160158 672
rect 166994 660 167000 672
rect 160152 632 167000 660
rect 160152 620 160158 632
rect 166994 620 167000 632
rect 167052 620 167058 672
rect 167178 620 167184 672
rect 167236 660 167242 672
rect 167236 632 169156 660
rect 167236 620 167242 632
rect 125226 592 125232 604
rect 116596 564 125232 592
rect 125226 552 125232 564
rect 125284 552 125290 604
rect 130562 552 130568 604
rect 130620 592 130626 604
rect 141786 592 141792 604
rect 130620 564 141792 592
rect 130620 552 130626 564
rect 141786 552 141792 564
rect 141844 552 141850 604
rect 142430 552 142436 604
rect 142488 592 142494 604
rect 150434 592 150440 604
rect 142488 564 150440 592
rect 142488 552 142494 564
rect 150434 552 150440 564
rect 150492 552 150498 604
rect 150618 552 150624 604
rect 150676 552 150682 604
rect 154206 552 154212 604
rect 154264 592 154270 604
rect 163866 592 163872 604
rect 154264 564 163872 592
rect 154264 552 154270 564
rect 163866 552 163872 564
rect 163924 552 163930 604
rect 120810 524 120816 536
rect 116504 496 120816 524
rect 120810 484 120816 496
rect 120868 484 120874 536
rect 124858 484 124864 536
rect 124916 524 124922 536
rect 136266 524 136272 536
rect 124916 496 136272 524
rect 124916 484 124922 496
rect 136266 484 136272 496
rect 136324 484 136330 536
rect 120074 416 120080 468
rect 120132 456 120138 468
rect 120132 428 127664 456
rect 120132 416 120138 428
rect 109126 348 109132 400
rect 109184 388 109190 400
rect 121914 388 121920 400
rect 109184 360 121920 388
rect 109184 348 109190 360
rect 121914 348 121920 360
rect 121972 348 121978 400
rect 122466 348 122472 400
rect 122524 388 122530 400
rect 127526 388 127532 400
rect 122524 360 127532 388
rect 122524 348 122530 360
rect 127526 348 127532 360
rect 127584 348 127590 400
rect 127636 388 127664 428
rect 131574 416 131580 468
rect 131632 456 131638 468
rect 142890 456 142896 468
rect 131632 428 142896 456
rect 131632 416 131638 428
rect 142890 416 142896 428
rect 142948 416 142954 468
rect 145742 416 145748 468
rect 145800 456 145806 468
rect 145800 428 150572 456
rect 145800 416 145806 428
rect 131942 388 131948 400
rect 127636 360 131948 388
rect 131942 348 131948 360
rect 132000 348 132006 400
rect 137462 348 137468 400
rect 137520 388 137526 400
rect 148502 388 148508 400
rect 137520 360 148508 388
rect 137520 348 137526 360
rect 148502 348 148508 360
rect 148560 348 148566 400
rect 106016 292 108988 320
rect 110690 280 110696 332
rect 110748 320 110754 332
rect 123018 320 123024 332
rect 110748 292 123024 320
rect 110748 280 110754 292
rect 123018 280 123024 292
rect 123076 280 123082 332
rect 125686 280 125692 332
rect 125744 320 125750 332
rect 137370 320 137376 332
rect 125744 292 137376 320
rect 125744 280 125750 292
rect 137370 280 137376 292
rect 137428 280 137434 332
rect 139026 280 139032 332
rect 139084 320 139090 332
rect 149330 320 149336 332
rect 139084 292 149336 320
rect 139084 280 139090 292
rect 149330 280 149336 292
rect 149388 280 149394 332
rect 28074 252 28080 264
rect 1544 224 19012 252
rect 21284 224 28080 252
rect 1544 212 1550 224
rect 3050 144 3056 196
rect 3108 184 3114 196
rect 18874 184 18880 196
rect 3108 156 18880 184
rect 3108 144 3114 156
rect 18874 144 18880 156
rect 18932 144 18938 196
rect 18984 184 19012 224
rect 28074 212 28080 224
rect 28132 212 28138 264
rect 44450 212 44456 264
rect 44508 252 44514 264
rect 61194 252 61200 264
rect 44508 224 61200 252
rect 44508 212 44514 224
rect 61194 212 61200 224
rect 61252 212 61258 264
rect 63402 212 63408 264
rect 63460 252 63466 264
rect 78858 252 78864 264
rect 63460 224 78864 252
rect 63460 212 63466 224
rect 78858 212 78864 224
rect 78916 212 78922 264
rect 81066 212 81072 264
rect 81124 252 81130 264
rect 94590 252 94596 264
rect 81124 224 94596 252
rect 81124 212 81130 224
rect 94590 212 94596 224
rect 94648 212 94654 264
rect 98454 212 98460 264
rect 98512 252 98518 264
rect 111978 252 111984 264
rect 98512 224 111984 252
rect 98512 212 98518 224
rect 111978 212 111984 224
rect 112036 212 112042 264
rect 114186 212 114192 264
rect 114244 252 114250 264
rect 126330 252 126336 264
rect 114244 224 126336 252
rect 114244 212 114250 224
rect 126330 212 126336 224
rect 126388 212 126394 264
rect 126790 212 126796 264
rect 126848 252 126854 264
rect 138474 252 138480 264
rect 126848 224 138480 252
rect 126848 212 126854 224
rect 138474 212 138480 224
rect 138532 212 138538 264
rect 21450 184 21456 196
rect 18984 156 21456 184
rect 21450 144 21456 156
rect 21508 144 21514 196
rect 27890 144 27896 196
rect 27948 184 27954 196
rect 45738 184 45744 196
rect 27948 156 45744 184
rect 27948 144 27954 156
rect 45738 144 45744 156
rect 45796 144 45802 196
rect 50338 144 50344 196
rect 50396 184 50402 196
rect 66530 184 66536 196
rect 50396 156 66536 184
rect 50396 144 50402 156
rect 66530 144 66536 156
rect 66588 144 66594 196
rect 68186 144 68192 196
rect 68244 184 68250 196
rect 83090 184 83096 196
rect 68244 156 83096 184
rect 68244 144 68250 156
rect 83090 144 83096 156
rect 83148 144 83154 196
rect 85850 144 85856 196
rect 85908 184 85914 196
rect 99650 184 99656 196
rect 85908 156 99656 184
rect 85908 144 85914 156
rect 99650 144 99656 156
rect 99708 144 99714 196
rect 102410 144 102416 196
rect 102468 184 102474 196
rect 115382 184 115388 196
rect 102468 156 115388 184
rect 102468 144 102474 156
rect 115382 144 115388 156
rect 115440 144 115446 196
rect 116578 144 116584 196
rect 116636 184 116642 196
rect 128538 184 128544 196
rect 116636 156 128544 184
rect 116636 144 116642 156
rect 128538 144 128544 156
rect 128596 144 128602 196
rect 133138 144 133144 196
rect 133196 184 133202 196
rect 143994 184 144000 196
rect 133196 156 144000 184
rect 133196 144 133202 156
rect 143994 144 144000 156
rect 144052 144 144058 196
rect 150544 184 150572 428
rect 150636 252 150664 552
rect 156414 416 156420 468
rect 156472 456 156478 468
rect 165890 456 165896 468
rect 156472 428 165896 456
rect 156472 416 156478 428
rect 165890 416 165896 428
rect 165948 416 165954 468
rect 155586 348 155592 400
rect 155644 388 155650 400
rect 165062 388 165068 400
rect 155644 360 165068 388
rect 155644 348 155650 360
rect 165062 348 165068 360
rect 165120 348 165126 400
rect 153194 280 153200 332
rect 153252 320 153258 332
rect 158714 320 158720 332
rect 153252 292 158720 320
rect 153252 280 153258 292
rect 158714 280 158720 292
rect 158772 280 158778 332
rect 159082 280 159088 332
rect 159140 320 159146 332
rect 168190 320 168196 332
rect 159140 292 168196 320
rect 159140 280 159146 292
rect 168190 280 168196 292
rect 168248 280 168254 332
rect 169128 320 169156 632
rect 169570 620 169576 672
rect 169628 660 169634 672
rect 175274 660 175280 672
rect 169628 632 175280 660
rect 169628 620 169634 632
rect 175274 620 175280 632
rect 175332 620 175338 672
rect 181714 660 181720 672
rect 175384 632 181720 660
rect 174262 552 174268 604
rect 174320 592 174326 604
rect 175384 592 175412 632
rect 181714 620 181720 632
rect 181772 620 181778 672
rect 182542 620 182548 672
rect 182600 660 182606 672
rect 187804 660 187832 700
rect 190362 688 190368 700
rect 190420 688 190426 740
rect 194410 688 194416 740
rect 194468 728 194474 740
rect 201402 728 201408 740
rect 194468 700 201408 728
rect 194468 688 194474 700
rect 201402 688 201408 700
rect 201460 688 201466 740
rect 201494 688 201500 740
rect 201552 728 201558 740
rect 205634 728 205640 740
rect 201552 700 205640 728
rect 201552 688 201558 700
rect 205634 688 205640 700
rect 205692 688 205698 740
rect 209774 688 209780 740
rect 209832 728 209838 740
rect 214834 728 214840 740
rect 209832 700 214840 728
rect 209832 688 209838 700
rect 214834 688 214840 700
rect 214892 688 214898 740
rect 215662 688 215668 740
rect 215720 728 215726 740
rect 220354 728 220360 740
rect 215720 700 220360 728
rect 215720 688 215726 700
rect 220354 688 220360 700
rect 220412 688 220418 740
rect 220446 688 220452 740
rect 220504 728 220510 740
rect 224770 728 224776 740
rect 220504 700 224776 728
rect 220504 688 220510 700
rect 224770 688 224776 700
rect 224828 688 224834 740
rect 233418 688 233424 740
rect 233476 728 233482 740
rect 237834 728 237840 740
rect 233476 700 237840 728
rect 233476 688 233482 700
rect 237834 688 237840 700
rect 237892 688 237898 740
rect 248782 688 248788 740
rect 248840 728 248846 740
rect 252186 728 252192 740
rect 248840 700 252192 728
rect 248840 688 248846 700
rect 252186 688 252192 700
rect 252244 688 252250 740
rect 318518 688 318524 740
rect 318576 728 318582 740
rect 319714 728 319720 740
rect 318576 700 319720 728
rect 318576 688 318582 700
rect 319714 688 319720 700
rect 319772 688 319778 740
rect 341702 688 341708 740
rect 341760 728 341766 740
rect 344554 728 344560 740
rect 341760 700 344560 728
rect 341760 688 341766 700
rect 344554 688 344560 700
rect 344612 688 344618 740
rect 350442 688 350448 740
rect 350500 728 350506 740
rect 354030 728 354036 740
rect 350500 700 354036 728
rect 350500 688 350506 700
rect 354030 688 354036 700
rect 354088 688 354094 740
rect 364886 688 364892 740
rect 364944 728 364950 740
rect 369394 728 369400 740
rect 364944 700 369400 728
rect 364944 688 364950 700
rect 369394 688 369400 700
rect 369452 688 369458 740
rect 380158 688 380164 740
rect 380216 728 380222 740
rect 384758 728 384764 740
rect 380216 700 384764 728
rect 380216 688 380222 700
rect 384758 688 384764 700
rect 384816 688 384822 740
rect 390646 688 390652 740
rect 390704 728 390710 740
rect 394234 728 394240 740
rect 390704 700 394240 728
rect 390704 688 390710 700
rect 394234 688 394240 700
rect 394292 688 394298 740
rect 396718 688 396724 740
rect 396776 728 396782 740
rect 400122 728 400128 740
rect 396776 700 400128 728
rect 396776 688 396782 700
rect 400122 688 400128 700
rect 400180 688 400186 740
rect 407758 688 407764 740
rect 407816 728 407822 740
rect 414290 728 414296 740
rect 407816 700 414296 728
rect 407816 688 407822 700
rect 414290 688 414296 700
rect 414348 688 414354 740
rect 414566 688 414572 740
rect 414624 728 414630 740
rect 422570 728 422576 740
rect 414624 700 422576 728
rect 414624 688 414630 700
rect 422570 688 422576 700
rect 422628 688 422634 740
rect 425422 688 425428 740
rect 425480 728 425486 740
rect 433242 728 433248 740
rect 425480 700 433248 728
rect 425480 688 425486 700
rect 433242 688 433248 700
rect 433300 688 433306 740
rect 448790 688 448796 740
rect 448848 728 448854 740
rect 459186 728 459192 740
rect 448848 700 459192 728
rect 448848 688 448854 700
rect 459186 688 459192 700
rect 459244 688 459250 740
rect 459830 688 459836 740
rect 459888 728 459894 740
rect 462976 728 463004 768
rect 471054 756 471060 768
rect 471112 756 471118 808
rect 481910 756 481916 808
rect 481968 796 481974 808
rect 494698 796 494704 808
rect 481968 768 494704 796
rect 481968 756 481974 768
rect 494698 756 494704 768
rect 494756 756 494762 808
rect 498470 756 498476 808
rect 498528 796 498534 808
rect 503622 796 503628 808
rect 498528 768 503628 796
rect 498528 756 498534 768
rect 503622 756 503628 768
rect 503680 756 503686 808
rect 459888 700 463004 728
rect 459888 688 459894 700
rect 463602 688 463608 740
rect 463660 728 463666 740
rect 463660 700 468708 728
rect 463660 688 463666 700
rect 182600 632 187832 660
rect 182600 620 182606 632
rect 188522 620 188528 672
rect 188580 660 188586 672
rect 188580 632 190454 660
rect 188580 620 188586 632
rect 174320 564 175412 592
rect 174320 552 174326 564
rect 176654 552 176660 604
rect 176712 592 176718 604
rect 184842 592 184848 604
rect 176712 564 184848 592
rect 176712 552 176718 564
rect 184842 552 184848 564
rect 184900 552 184906 604
rect 189718 552 189724 604
rect 189776 552 189782 604
rect 190426 592 190454 632
rect 195606 620 195612 672
rect 195664 660 195670 672
rect 202506 660 202512 672
rect 195664 632 202512 660
rect 195664 620 195670 632
rect 202506 620 202512 632
rect 202564 620 202570 672
rect 204254 660 204260 672
rect 202616 632 204260 660
rect 195882 592 195888 604
rect 190426 564 195888 592
rect 195882 552 195888 564
rect 195940 552 195946 604
rect 200298 552 200304 604
rect 200356 592 200362 604
rect 202616 592 202644 632
rect 204254 620 204260 632
rect 204312 620 204318 672
rect 207382 620 207388 672
rect 207440 660 207446 672
rect 211614 660 211620 672
rect 207440 632 211620 660
rect 207440 620 207446 632
rect 211614 620 211620 632
rect 211672 620 211678 672
rect 212166 620 212172 672
rect 212224 660 212230 672
rect 215294 660 215300 672
rect 212224 632 215300 660
rect 212224 620 212230 632
rect 215294 620 215300 632
rect 215352 620 215358 672
rect 216858 620 216864 672
rect 216916 660 216922 672
rect 221458 660 221464 672
rect 216916 632 221464 660
rect 216916 620 216922 632
rect 221458 620 221464 632
rect 221516 620 221522 672
rect 226334 620 226340 672
rect 226392 660 226398 672
rect 231210 660 231216 672
rect 226392 632 231216 660
rect 226392 620 226398 632
rect 231210 620 231216 632
rect 231268 620 231274 672
rect 234614 620 234620 672
rect 234672 660 234678 672
rect 238938 660 238944 672
rect 234672 632 238944 660
rect 234672 620 234678 632
rect 238938 620 238944 632
rect 238996 620 239002 672
rect 240502 620 240508 672
rect 240560 660 240566 672
rect 244458 660 244464 672
rect 240560 632 244464 660
rect 240560 620 240566 632
rect 244458 620 244464 632
rect 244516 620 244522 672
rect 245194 620 245200 672
rect 245252 660 245258 672
rect 248874 660 248880 672
rect 245252 632 248880 660
rect 245252 620 245258 632
rect 248874 620 248880 632
rect 248932 620 248938 672
rect 262950 620 262956 672
rect 263008 660 263014 672
rect 265434 660 265440 672
rect 263008 632 265440 660
rect 263008 620 263014 632
rect 265434 620 265440 632
rect 265492 620 265498 672
rect 333974 620 333980 672
rect 334032 660 334038 672
rect 336274 660 336280 672
rect 334032 632 336280 660
rect 334032 620 334038 632
rect 336274 620 336280 632
rect 336332 620 336338 672
rect 339494 620 339500 672
rect 339552 660 339558 672
rect 342162 660 342168 672
rect 339552 632 342168 660
rect 339552 620 339558 632
rect 342162 620 342168 632
rect 342220 620 342226 672
rect 349890 620 349896 672
rect 349948 660 349954 672
rect 351638 660 351644 672
rect 349948 632 351644 660
rect 349948 620 349954 632
rect 351638 620 351644 632
rect 351696 620 351702 672
rect 360470 620 360476 672
rect 360528 660 360534 672
rect 364610 660 364616 672
rect 360528 632 364616 660
rect 360528 620 360534 632
rect 364610 620 364616 632
rect 364668 620 364674 672
rect 366174 620 366180 672
rect 366232 660 366238 672
rect 368198 660 368204 672
rect 366232 632 368204 660
rect 366232 620 366238 632
rect 368198 620 368204 632
rect 368256 620 368262 672
rect 368290 620 368296 672
rect 368348 660 368354 672
rect 372890 660 372896 672
rect 368348 632 372896 660
rect 368348 620 368354 632
rect 372890 620 372896 632
rect 372948 620 372954 672
rect 378502 620 378508 672
rect 378560 660 378566 672
rect 381170 660 381176 672
rect 378560 632 381176 660
rect 378560 620 378566 632
rect 381170 620 381176 632
rect 381228 620 381234 672
rect 384666 620 384672 672
rect 384724 660 384730 672
rect 384724 632 389036 660
rect 384724 620 384730 632
rect 200356 564 202644 592
rect 200356 552 200362 564
rect 202690 552 202696 604
rect 202748 592 202754 604
rect 209130 592 209136 604
rect 202748 564 209136 592
rect 202748 552 202754 564
rect 209130 552 209136 564
rect 209188 552 209194 604
rect 213362 552 213368 604
rect 213420 592 213426 604
rect 216674 592 216680 604
rect 213420 564 216680 592
rect 213420 552 213426 564
rect 216674 552 216680 564
rect 216732 552 216738 604
rect 218054 552 218060 604
rect 218112 552 218118 604
rect 221550 552 221556 604
rect 221608 592 221614 604
rect 224954 592 224960 604
rect 221608 564 224960 592
rect 221608 552 221614 564
rect 224954 552 224960 564
rect 225012 552 225018 604
rect 227530 552 227536 604
rect 227588 592 227594 604
rect 230566 592 230572 604
rect 227588 564 230572 592
rect 227588 552 227594 564
rect 230566 552 230572 564
rect 230624 552 230630 604
rect 232222 552 232228 604
rect 232280 592 232286 604
rect 234706 592 234712 604
rect 232280 564 234712 592
rect 232280 552 232286 564
rect 234706 552 234712 564
rect 234764 552 234770 604
rect 237006 552 237012 604
rect 237064 592 237070 604
rect 241146 592 241152 604
rect 237064 564 241152 592
rect 237064 552 237070 564
rect 241146 552 241152 564
rect 241204 552 241210 604
rect 241698 552 241704 604
rect 241756 592 241762 604
rect 245562 592 245568 604
rect 241756 564 245568 592
rect 241756 552 241762 564
rect 245562 552 245568 564
rect 245620 552 245626 604
rect 246390 552 246396 604
rect 246448 592 246454 604
rect 250070 592 250076 604
rect 246448 564 250076 592
rect 246448 552 246454 564
rect 250070 552 250076 564
rect 250128 552 250134 604
rect 251174 552 251180 604
rect 251232 592 251238 604
rect 254394 592 254400 604
rect 251232 564 254400 592
rect 251232 552 251238 564
rect 254394 552 254400 564
rect 254452 552 254458 604
rect 254670 552 254676 604
rect 254728 592 254734 604
rect 257706 592 257712 604
rect 254728 564 257712 592
rect 254728 552 254734 564
rect 257706 552 257712 564
rect 257764 552 257770 604
rect 258258 552 258264 604
rect 258316 592 258322 604
rect 261018 592 261024 604
rect 258316 564 261024 592
rect 258316 552 258322 564
rect 261018 552 261024 564
rect 261076 552 261082 604
rect 264146 552 264152 604
rect 264204 592 264210 604
rect 266630 592 266636 604
rect 264204 564 266636 592
rect 264204 552 264210 564
rect 266630 552 266636 564
rect 266688 552 266694 604
rect 268838 552 268844 604
rect 268896 592 268902 604
rect 270954 592 270960 604
rect 268896 564 270960 592
rect 268896 552 268902 564
rect 270954 552 270960 564
rect 271012 552 271018 604
rect 277118 552 277124 604
rect 277176 592 277182 604
rect 278682 592 278688 604
rect 277176 564 278688 592
rect 277176 552 277182 564
rect 278682 552 278688 564
rect 278740 552 278746 604
rect 307478 552 307484 604
rect 307536 592 307542 604
rect 307938 592 307944 604
rect 307536 564 307944 592
rect 307536 552 307542 564
rect 307938 552 307944 564
rect 307996 552 308002 604
rect 312998 552 313004 604
rect 313056 592 313062 604
rect 313826 592 313832 604
rect 313056 564 313832 592
rect 313056 552 313062 564
rect 313826 552 313832 564
rect 313884 552 313890 604
rect 315206 552 315212 604
rect 315264 592 315270 604
rect 316218 592 316224 604
rect 315264 564 316224 592
rect 315264 552 315270 564
rect 316218 552 316224 564
rect 316276 552 316282 604
rect 317230 552 317236 604
rect 317288 592 317294 604
rect 318518 592 318524 604
rect 317288 564 318524 592
rect 317288 552 317294 564
rect 318518 552 318524 564
rect 318576 552 318582 604
rect 319622 552 319628 604
rect 319680 592 319686 604
rect 320910 592 320916 604
rect 319680 564 320916 592
rect 319680 552 319686 564
rect 320910 552 320916 564
rect 320968 552 320974 604
rect 324038 552 324044 604
rect 324096 592 324102 604
rect 325602 592 325608 604
rect 324096 564 325608 592
rect 324096 552 324102 564
rect 325602 552 325608 564
rect 325660 552 325666 604
rect 326246 552 326252 604
rect 326304 592 326310 604
rect 327994 592 328000 604
rect 326304 564 328000 592
rect 326304 552 326310 564
rect 327994 552 328000 564
rect 328052 552 328058 604
rect 328362 552 328368 604
rect 328420 592 328426 604
rect 330386 592 330392 604
rect 328420 564 330392 592
rect 328420 552 328426 564
rect 330386 552 330392 564
rect 330444 552 330450 604
rect 332870 552 332876 604
rect 332928 592 332934 604
rect 335078 592 335084 604
rect 332928 564 335084 592
rect 332928 552 332934 564
rect 335078 552 335084 564
rect 335136 552 335142 604
rect 337286 552 337292 604
rect 337344 592 337350 604
rect 339862 592 339868 604
rect 337344 564 339868 592
rect 337344 552 337350 564
rect 339862 552 339868 564
rect 339920 552 339926 604
rect 343910 552 343916 604
rect 343968 592 343974 604
rect 346946 592 346952 604
rect 343968 564 346952 592
rect 343968 552 343974 564
rect 346946 552 346952 564
rect 347004 552 347010 604
rect 348786 552 348792 604
rect 348844 592 348850 604
rect 350442 592 350448 604
rect 348844 564 350448 592
rect 348844 552 348850 564
rect 350442 552 350448 564
rect 350500 552 350506 604
rect 355778 552 355784 604
rect 355836 592 355842 604
rect 356330 592 356336 604
rect 355836 564 356336 592
rect 355836 552 355842 564
rect 356330 552 356336 564
rect 356388 552 356394 604
rect 357158 552 357164 604
rect 357216 592 357222 604
rect 361114 592 361120 604
rect 357216 564 361120 592
rect 357216 552 357222 564
rect 361114 552 361120 564
rect 361172 552 361178 604
rect 363506 552 363512 604
rect 363564 592 363570 604
rect 367002 592 367008 604
rect 363564 564 367008 592
rect 363564 552 363570 564
rect 367002 552 367008 564
rect 367060 552 367066 604
rect 369762 552 369768 604
rect 369820 592 369826 604
rect 370590 592 370596 604
rect 369820 564 370596 592
rect 369820 552 369826 564
rect 370590 552 370596 564
rect 370648 552 370654 604
rect 372706 552 372712 604
rect 372764 592 372770 604
rect 375282 592 375288 604
rect 372764 564 375288 592
rect 372764 552 372770 564
rect 375282 552 375288 564
rect 375340 552 375346 604
rect 376662 552 376668 604
rect 376720 592 376726 604
rect 379974 592 379980 604
rect 376720 564 379980 592
rect 376720 552 376726 564
rect 379974 552 379980 564
rect 380032 552 380038 604
rect 382274 552 382280 604
rect 382332 592 382338 604
rect 385954 592 385960 604
rect 382332 564 385960 592
rect 382332 552 382338 564
rect 385954 552 385960 564
rect 386012 552 386018 604
rect 389008 592 389036 632
rect 389082 620 389088 672
rect 389140 660 389146 672
rect 395338 660 395344 672
rect 389140 632 395344 660
rect 389140 620 389146 632
rect 395338 620 395344 632
rect 395396 620 395402 672
rect 395798 620 395804 672
rect 395856 660 395862 672
rect 395856 632 398696 660
rect 395856 620 395862 632
rect 390646 592 390652 604
rect 389008 564 390652 592
rect 390646 552 390652 564
rect 390704 552 390710 604
rect 394418 552 394424 604
rect 394476 592 394482 604
rect 397730 592 397736 604
rect 394476 564 397736 592
rect 394476 552 394482 564
rect 397730 552 397736 564
rect 397788 552 397794 604
rect 398668 592 398696 632
rect 398742 620 398748 672
rect 398800 660 398806 672
rect 403618 660 403624 672
rect 398800 632 403624 660
rect 398800 620 398806 632
rect 403618 620 403624 632
rect 403676 620 403682 672
rect 407022 620 407028 672
rect 407080 660 407086 672
rect 410794 660 410800 672
rect 407080 632 410800 660
rect 407080 620 407086 632
rect 410794 620 410800 632
rect 410852 620 410858 672
rect 417786 620 417792 672
rect 417844 660 417850 672
rect 417844 632 419120 660
rect 417844 620 417850 632
rect 402514 592 402520 604
rect 398668 564 402520 592
rect 402514 552 402520 564
rect 402572 552 402578 604
rect 406010 552 406016 604
rect 406068 552 406074 604
rect 409782 552 409788 604
rect 409840 592 409846 604
rect 415486 592 415492 604
rect 409840 564 415492 592
rect 409840 552 409846 564
rect 415486 552 415492 564
rect 415544 552 415550 604
rect 417878 552 417884 604
rect 417936 552 417942 604
rect 178034 484 178040 536
rect 178092 524 178098 536
rect 185946 524 185952 536
rect 178092 496 185952 524
rect 178092 484 178098 496
rect 185946 484 185952 496
rect 186004 484 186010 536
rect 189736 524 189764 552
rect 196986 524 196992 536
rect 189736 496 196992 524
rect 196986 484 196992 496
rect 197044 484 197050 536
rect 172146 416 172152 468
rect 172204 456 172210 468
rect 180426 456 180432 468
rect 172204 428 180432 456
rect 172204 416 172210 428
rect 180426 416 180432 428
rect 180484 416 180490 468
rect 192202 416 192208 468
rect 192260 456 192266 468
rect 199286 456 199292 468
rect 192260 428 199292 456
rect 192260 416 192266 428
rect 199286 416 199292 428
rect 199344 416 199350 468
rect 170582 348 170588 400
rect 170640 388 170646 400
rect 179322 388 179328 400
rect 170640 360 179328 388
rect 170640 348 170646 360
rect 179322 348 179328 360
rect 179380 348 179386 400
rect 196986 348 196992 400
rect 197044 388 197050 400
rect 203610 388 203616 400
rect 197044 360 203616 388
rect 197044 348 197050 360
rect 203610 348 203616 360
rect 203668 348 203674 400
rect 208762 348 208768 400
rect 208820 388 208826 400
rect 213730 388 213736 400
rect 208820 360 213736 388
rect 208820 348 208826 360
rect 213730 348 213736 360
rect 213788 348 213794 400
rect 176010 320 176016 332
rect 169128 292 176016 320
rect 176010 280 176016 292
rect 176068 280 176074 332
rect 178862 280 178868 332
rect 178920 320 178926 332
rect 187050 320 187056 332
rect 178920 292 187056 320
rect 178920 280 178926 292
rect 187050 280 187056 292
rect 187108 280 187114 332
rect 205266 280 205272 332
rect 205324 320 205330 332
rect 211338 320 211344 332
rect 205324 292 211344 320
rect 205324 280 205330 292
rect 211338 280 211344 292
rect 211396 280 211402 332
rect 160554 252 160560 264
rect 150636 224 160560 252
rect 160554 212 160560 224
rect 160612 212 160618 264
rect 162302 212 162308 264
rect 162360 252 162366 264
rect 171594 252 171600 264
rect 162360 224 171600 252
rect 162360 212 162366 224
rect 171594 212 171600 224
rect 171652 212 171658 264
rect 186314 212 186320 264
rect 186372 252 186378 264
rect 193674 252 193680 264
rect 186372 224 193680 252
rect 186372 212 186378 224
rect 193674 212 193680 224
rect 193732 212 193738 264
rect 198090 212 198096 264
rect 198148 252 198154 264
rect 204714 252 204720 264
rect 198148 224 204720 252
rect 198148 212 198154 224
rect 204714 212 204720 224
rect 204772 212 204778 264
rect 206370 212 206376 264
rect 206428 252 206434 264
rect 212442 252 212448 264
rect 206428 224 212448 252
rect 206428 212 206434 224
rect 212442 212 212448 224
rect 212500 212 212506 264
rect 156138 184 156144 196
rect 150544 156 156144 184
rect 156138 144 156144 156
rect 156196 144 156202 196
rect 163866 144 163872 196
rect 163924 184 163930 196
rect 172698 184 172704 196
rect 163924 156 172704 184
rect 163924 144 163930 156
rect 172698 144 172704 156
rect 172756 144 172762 196
rect 175642 144 175648 196
rect 175700 184 175706 196
rect 183554 184 183560 196
rect 175700 156 183560 184
rect 175700 144 175706 156
rect 183554 144 183560 156
rect 183612 144 183618 196
rect 187142 144 187148 196
rect 187200 184 187206 196
rect 194778 184 194784 196
rect 187200 156 194784 184
rect 187200 144 187206 156
rect 194778 144 194784 156
rect 194836 144 194842 196
rect 198918 144 198924 196
rect 198976 184 198982 196
rect 205818 184 205824 196
rect 198976 156 205824 184
rect 198976 144 198982 156
rect 205818 144 205824 156
rect 205876 144 205882 196
rect 218072 184 218100 552
rect 401594 484 401600 536
rect 401652 524 401658 536
rect 406028 524 406056 552
rect 401652 496 406056 524
rect 401652 484 401658 496
rect 225322 416 225328 468
rect 225380 456 225386 468
rect 230106 456 230112 468
rect 225380 428 230112 456
rect 225380 416 225386 428
rect 230106 416 230112 428
rect 230164 416 230170 468
rect 239490 416 239496 468
rect 239548 456 239554 468
rect 243354 456 243360 468
rect 239548 428 243360 456
rect 239548 416 239554 428
rect 243354 416 243360 428
rect 243412 416 243418 468
rect 361482 416 361488 468
rect 361540 456 361546 468
rect 365622 456 365628 468
rect 361540 428 365628 456
rect 361540 416 361546 428
rect 365622 416 365628 428
rect 365680 416 365686 468
rect 371510 416 371516 468
rect 371568 456 371574 468
rect 376294 456 376300 468
rect 371568 428 376300 456
rect 371568 416 371574 428
rect 376294 416 376300 428
rect 376352 416 376358 468
rect 377030 416 377036 468
rect 377088 456 377094 468
rect 382182 456 382188 468
rect 377088 428 382188 456
rect 377088 416 377094 428
rect 382182 416 382188 428
rect 382240 416 382246 468
rect 387886 416 387892 468
rect 387944 456 387950 468
rect 392854 456 392860 468
rect 387944 428 392860 456
rect 387944 416 387950 428
rect 392854 416 392860 428
rect 392912 416 392918 468
rect 219434 348 219440 400
rect 219492 388 219498 400
rect 222562 388 222568 400
rect 219492 360 222568 388
rect 219492 348 219498 360
rect 222562 348 222568 360
rect 222620 348 222626 400
rect 222930 348 222936 400
rect 222988 388 222994 400
rect 226518 388 226524 400
rect 222988 360 226524 388
rect 222988 348 222994 360
rect 226518 348 226524 360
rect 226576 348 226582 400
rect 231210 348 231216 400
rect 231268 388 231274 400
rect 235626 388 235632 400
rect 231268 360 235632 388
rect 231268 348 231274 360
rect 235626 348 235632 360
rect 235684 348 235690 400
rect 235994 348 236000 400
rect 236052 388 236058 400
rect 240042 388 240048 400
rect 236052 360 240048 388
rect 236052 348 236058 360
rect 240042 348 240048 360
rect 240100 348 240106 400
rect 244274 348 244280 400
rect 244332 388 244338 400
rect 247770 388 247776 400
rect 244332 360 247776 388
rect 244332 348 244338 360
rect 247770 348 247776 360
rect 247828 348 247834 400
rect 252554 348 252560 400
rect 252612 388 252618 400
rect 255498 388 255504 400
rect 252612 360 255504 388
rect 252612 348 252618 360
rect 255498 348 255504 360
rect 255556 348 255562 400
rect 256050 348 256056 400
rect 256108 388 256114 400
rect 258810 388 258816 400
rect 256108 360 258816 388
rect 256108 348 256114 360
rect 258810 348 258816 360
rect 258868 348 258874 400
rect 260834 348 260840 400
rect 260892 388 260898 400
rect 263226 388 263232 400
rect 260892 360 263232 388
rect 260892 348 260898 360
rect 263226 348 263232 360
rect 263284 348 263290 400
rect 270218 348 270224 400
rect 270276 388 270282 400
rect 272058 388 272064 400
rect 270276 360 272064 388
rect 270276 348 270282 360
rect 272058 348 272064 360
rect 272116 348 272122 400
rect 311802 348 311808 400
rect 311860 388 311866 400
rect 312446 388 312452 400
rect 311860 360 312452 388
rect 311860 348 311866 360
rect 312446 348 312452 360
rect 312504 348 312510 400
rect 314102 348 314108 400
rect 314160 388 314166 400
rect 314838 388 314844 400
rect 314160 360 314844 388
rect 314160 348 314166 360
rect 314838 348 314844 360
rect 314896 348 314902 400
rect 321830 348 321836 400
rect 321888 388 321894 400
rect 323118 388 323124 400
rect 321888 360 323124 388
rect 321888 348 321894 360
rect 323118 348 323124 360
rect 323176 348 323182 400
rect 327350 348 327356 400
rect 327408 388 327414 400
rect 329006 388 329012 400
rect 327408 360 329012 388
rect 327408 348 327414 360
rect 329006 348 329012 360
rect 329064 348 329070 400
rect 330662 348 330668 400
rect 330720 388 330726 400
rect 332502 388 332508 400
rect 330720 360 332508 388
rect 330720 348 330726 360
rect 332502 348 332508 360
rect 332560 348 332566 400
rect 336458 348 336464 400
rect 336516 388 336522 400
rect 337286 388 337292 400
rect 336516 360 337292 388
rect 336516 348 336522 360
rect 337286 348 337292 360
rect 337344 348 337350 400
rect 338390 348 338396 400
rect 338448 388 338454 400
rect 340782 388 340788 400
rect 338448 360 340788 388
rect 338448 348 338454 360
rect 340782 348 340788 360
rect 340840 348 340846 400
rect 347590 348 347596 400
rect 347648 388 347654 400
rect 349062 388 349068 400
rect 347648 360 349068 388
rect 347648 348 347654 360
rect 349062 348 349068 360
rect 349120 348 349126 400
rect 355870 348 355876 400
rect 355928 388 355934 400
rect 359734 388 359740 400
rect 355928 360 359740 388
rect 355928 348 355934 360
rect 359734 348 359740 360
rect 359792 348 359798 400
rect 360102 348 360108 400
rect 360160 388 360166 400
rect 362126 388 362132 400
rect 360160 360 362132 388
rect 360160 348 360166 360
rect 362126 348 362132 360
rect 362184 348 362190 400
rect 362494 348 362500 400
rect 362552 388 362558 400
rect 363690 388 363696 400
rect 362552 360 363696 388
rect 362552 348 362558 360
rect 363690 348 363696 360
rect 363748 348 363754 400
rect 370222 348 370228 400
rect 370280 388 370286 400
rect 373902 388 373908 400
rect 370280 360 373908 388
rect 370280 348 370286 360
rect 373902 348 373908 360
rect 373960 348 373966 400
rect 375098 348 375104 400
rect 375156 388 375162 400
rect 378686 388 378692 400
rect 375156 360 378692 388
rect 375156 348 375162 360
rect 378686 348 378692 360
rect 378744 348 378750 400
rect 392486 348 392492 400
rect 392544 388 392550 400
rect 398742 388 398748 400
rect 392544 360 398748 388
rect 392544 348 392550 360
rect 398742 348 398748 360
rect 398800 348 398806 400
rect 399846 348 399852 400
rect 399904 388 399910 400
rect 404630 388 404636 400
rect 399904 360 404636 388
rect 399904 348 399910 360
rect 404630 348 404636 360
rect 404688 348 404694 400
rect 404262 280 404268 332
rect 404320 320 404326 332
rect 409414 320 409420 332
rect 404320 292 409420 320
rect 404320 280 404326 292
rect 409414 280 409420 292
rect 409472 280 409478 332
rect 410150 280 410156 332
rect 410208 320 410214 332
rect 417896 320 417924 552
rect 410208 292 417924 320
rect 419092 320 419120 632
rect 428734 620 428740 672
rect 428792 660 428798 672
rect 434438 660 434444 672
rect 428792 632 434444 660
rect 428792 620 428798 632
rect 434438 620 434444 632
rect 434496 620 434502 672
rect 437934 660 437940 672
rect 435376 632 437940 660
rect 421190 552 421196 604
rect 421248 592 421254 604
rect 429654 592 429660 604
rect 421248 564 429660 592
rect 421248 552 421254 564
rect 429654 552 429660 564
rect 429712 552 429718 604
rect 435376 592 435404 632
rect 437934 620 437940 632
rect 437992 620 437998 672
rect 438946 620 438952 672
rect 439004 660 439010 672
rect 441522 660 441528 672
rect 439004 632 441528 660
rect 439004 620 439010 632
rect 441522 620 441528 632
rect 441580 620 441586 672
rect 442902 620 442908 672
rect 442960 660 442966 672
rect 442960 632 447640 660
rect 442960 620 442966 632
rect 435542 592 435548 604
rect 431926 564 435404 592
rect 419994 416 420000 468
rect 420052 456 420058 468
rect 428642 456 428648 468
rect 420052 428 428648 456
rect 420052 416 420058 428
rect 428642 416 428648 428
rect 428700 416 428706 468
rect 429838 416 429844 468
rect 429896 456 429902 468
rect 431926 456 431954 564
rect 429896 428 431954 456
rect 435514 552 435548 592
rect 435600 552 435606 604
rect 437750 552 437756 604
rect 437808 592 437814 604
rect 447410 592 447416 604
rect 437808 564 447416 592
rect 437808 552 437814 564
rect 447410 552 447416 564
rect 447468 552 447474 604
rect 447612 592 447640 632
rect 447686 620 447692 672
rect 447744 660 447750 672
rect 458082 660 458088 672
rect 447744 632 458088 660
rect 447744 620 447750 632
rect 458082 620 458088 632
rect 458140 620 458146 672
rect 458726 620 458732 672
rect 458784 660 458790 672
rect 467282 660 467288 672
rect 458784 632 467288 660
rect 458784 620 458790 632
rect 467282 620 467288 632
rect 467340 620 467346 672
rect 468570 660 468576 672
rect 467392 632 468576 660
rect 449802 592 449808 604
rect 447612 564 449808 592
rect 449802 552 449808 564
rect 449860 552 449866 604
rect 450906 552 450912 604
rect 450964 552 450970 604
rect 451182 552 451188 604
rect 451240 592 451246 604
rect 452102 592 452108 604
rect 451240 564 452108 592
rect 451240 552 451246 564
rect 452102 552 452108 564
rect 452160 552 452166 604
rect 452562 552 452568 604
rect 452620 592 452626 604
rect 461578 592 461584 604
rect 452620 564 461584 592
rect 452620 552 452626 564
rect 461578 552 461584 564
rect 461636 552 461642 604
rect 429896 416 429902 428
rect 419166 348 419172 400
rect 419224 388 419230 400
rect 427078 388 427084 400
rect 419224 360 427084 388
rect 419224 348 419230 360
rect 427078 348 427084 360
rect 427136 348 427142 400
rect 435514 388 435542 552
rect 436554 484 436560 536
rect 436612 524 436618 536
rect 446030 524 446036 536
rect 436612 496 446036 524
rect 436612 484 436618 496
rect 446030 484 446036 496
rect 446088 484 446094 536
rect 450924 456 450952 552
rect 454310 484 454316 536
rect 454368 524 454374 536
rect 464982 524 464988 536
rect 454368 496 464988 524
rect 454368 484 454374 496
rect 464982 484 464988 496
rect 465040 484 465046 536
rect 446232 428 450952 456
rect 429488 360 435542 388
rect 425974 320 425980 332
rect 419092 292 425980 320
rect 410208 280 410214 292
rect 425974 280 425980 292
rect 426032 280 426038 332
rect 426710 280 426716 332
rect 426768 320 426774 332
rect 429488 320 429516 360
rect 435726 348 435732 400
rect 435784 388 435790 400
rect 445202 388 445208 400
rect 435784 360 445208 388
rect 435784 348 435790 360
rect 445202 348 445208 360
rect 445260 348 445266 400
rect 426768 292 429516 320
rect 426768 280 426774 292
rect 431126 280 431132 332
rect 431184 320 431190 332
rect 440142 320 440148 332
rect 431184 292 440148 320
rect 431184 280 431190 292
rect 440142 280 440148 292
rect 440200 280 440206 332
rect 441062 280 441068 332
rect 441120 320 441126 332
rect 446232 320 446260 428
rect 451090 416 451096 468
rect 451148 456 451154 468
rect 453482 456 453488 468
rect 451148 428 453488 456
rect 451148 416 451154 428
rect 453482 416 453488 428
rect 453540 416 453546 468
rect 457622 416 457628 468
rect 457680 456 457686 468
rect 467392 456 467420 632
rect 468570 620 468576 632
rect 468628 620 468634 672
rect 467466 552 467472 604
rect 467524 552 467530 604
rect 468680 592 468708 700
rect 480806 688 480812 740
rect 480864 728 480870 740
rect 493502 728 493508 740
rect 480864 700 493508 728
rect 480864 688 480870 700
rect 493502 688 493508 700
rect 493560 688 493566 740
rect 499390 728 499396 740
rect 497292 700 499396 728
rect 469766 620 469772 672
rect 469824 660 469830 672
rect 481726 660 481732 672
rect 469824 632 481732 660
rect 469824 620 469830 632
rect 481726 620 481732 632
rect 481784 620 481790 672
rect 482922 620 482928 672
rect 482980 660 482986 672
rect 485498 660 485504 672
rect 482980 632 485504 660
rect 482980 620 482986 632
rect 485498 620 485504 632
rect 485556 620 485562 672
rect 485746 632 486280 660
rect 473446 592 473452 604
rect 468680 564 473452 592
rect 473446 552 473452 564
rect 473504 552 473510 604
rect 474182 552 474188 604
rect 474240 592 474246 604
rect 485746 592 485774 632
rect 474240 564 485774 592
rect 486252 592 486280 632
rect 486326 620 486332 672
rect 486384 660 486390 672
rect 497292 660 497320 700
rect 499390 688 499396 700
rect 499448 688 499454 740
rect 503732 728 503760 836
rect 504174 824 504180 836
rect 504232 824 504238 876
rect 507302 824 507308 876
rect 507360 864 507366 876
rect 521838 864 521844 876
rect 507360 836 521844 864
rect 507360 824 507366 836
rect 521838 824 521844 836
rect 521896 824 521902 876
rect 531590 824 531596 876
rect 531648 864 531654 876
rect 547874 864 547880 876
rect 531648 836 547880 864
rect 531648 824 531654 836
rect 547874 824 547880 836
rect 547932 824 547938 876
rect 552566 824 552572 876
rect 552624 864 552630 876
rect 570322 864 570328 876
rect 552624 836 570328 864
rect 552624 824 552630 836
rect 570322 824 570328 836
rect 570380 824 570386 876
rect 503898 756 503904 808
rect 503956 796 503962 808
rect 512454 796 512460 808
rect 503956 768 512460 796
rect 503956 756 503962 768
rect 512454 756 512460 768
rect 512512 756 512518 808
rect 517238 756 517244 808
rect 517296 796 517302 808
rect 532326 796 532332 808
rect 517296 768 532332 796
rect 517296 756 517302 768
rect 532326 756 532332 768
rect 532384 756 532390 808
rect 532528 768 538214 796
rect 506474 728 506480 740
rect 503732 700 506480 728
rect 506474 688 506480 700
rect 506532 688 506538 740
rect 515030 688 515036 740
rect 515088 728 515094 740
rect 530118 728 530124 740
rect 515088 700 530124 728
rect 515088 688 515094 700
rect 530118 688 530124 700
rect 530176 688 530182 740
rect 530486 688 530492 740
rect 530544 728 530550 740
rect 532528 728 532556 768
rect 530544 700 532556 728
rect 530544 688 530550 700
rect 532602 688 532608 740
rect 532660 728 532666 740
rect 538186 728 538214 768
rect 542630 756 542636 808
rect 542688 796 542694 808
rect 559098 796 559104 808
rect 542688 768 559104 796
rect 542688 756 542694 768
rect 559098 756 559104 768
rect 559156 756 559162 808
rect 559190 756 559196 808
rect 559248 796 559254 808
rect 577406 796 577412 808
rect 559248 768 577412 796
rect 559248 756 559254 768
rect 577406 756 577412 768
rect 577464 756 577470 808
rect 546678 728 546684 740
rect 532660 700 535500 728
rect 538186 700 546684 728
rect 532660 688 532666 700
rect 486384 632 497320 660
rect 486384 620 486390 632
rect 497366 620 497372 672
rect 497424 660 497430 672
rect 511258 660 511264 672
rect 497424 632 511264 660
rect 497424 620 497430 632
rect 511258 620 511264 632
rect 511316 620 511322 672
rect 513926 620 513932 672
rect 513984 660 513990 672
rect 513984 632 518894 660
rect 513984 620 513990 632
rect 486418 592 486424 604
rect 486252 564 486424 592
rect 474240 552 474246 564
rect 486418 552 486424 564
rect 486476 552 486482 604
rect 489638 552 489644 604
rect 489696 592 489702 604
rect 502978 592 502984 604
rect 489696 564 502984 592
rect 489696 552 489702 564
rect 502978 552 502984 564
rect 503036 552 503042 604
rect 517146 592 517152 604
rect 506032 564 517152 592
rect 457680 428 467420 456
rect 457680 416 457686 428
rect 446582 348 446588 400
rect 446640 388 446646 400
rect 456702 388 456708 400
rect 446640 360 456708 388
rect 446640 348 446646 360
rect 456702 348 456708 360
rect 456760 348 456766 400
rect 441120 292 446260 320
rect 441120 280 441126 292
rect 453114 280 453120 332
rect 453172 320 453178 332
rect 464154 320 464160 332
rect 453172 292 464160 320
rect 453172 280 453178 292
rect 464154 280 464160 292
rect 464212 280 464218 332
rect 237926 212 237932 264
rect 237984 252 237990 264
rect 242250 252 242256 264
rect 237984 224 242256 252
rect 237984 212 237990 224
rect 242250 212 242256 224
rect 242308 212 242314 264
rect 353846 212 353852 264
rect 353904 252 353910 264
rect 357342 252 357348 264
rect 353904 224 357348 252
rect 353904 212 353910 224
rect 357342 212 357348 224
rect 357400 212 357406 264
rect 390278 212 390284 264
rect 390336 252 390342 264
rect 396350 252 396356 264
rect 390336 224 396356 252
rect 390336 212 390342 224
rect 396350 212 396356 224
rect 396408 212 396414 264
rect 401502 212 401508 264
rect 401560 252 401566 264
rect 408586 252 408592 264
rect 401560 224 408592 252
rect 401560 212 401566 224
rect 408586 212 408592 224
rect 408644 212 408650 264
rect 412358 212 412364 264
rect 412416 252 412422 264
rect 420362 252 420368 264
rect 412416 224 420368 252
rect 412416 212 412422 224
rect 420362 212 420368 224
rect 420420 212 420426 264
rect 423398 212 423404 264
rect 423456 252 423462 264
rect 431862 252 431868 264
rect 423456 224 431868 252
rect 423456 212 423462 224
rect 431862 212 431868 224
rect 431920 212 431926 264
rect 434622 212 434628 264
rect 434680 252 434686 264
rect 443638 252 443644 264
rect 434680 224 443644 252
rect 434680 212 434686 224
rect 443638 212 443644 224
rect 443696 212 443702 264
rect 445478 212 445484 264
rect 445536 252 445542 264
rect 455874 252 455880 264
rect 445536 224 455880 252
rect 445536 212 445542 224
rect 455874 212 455880 224
rect 455932 212 455938 264
rect 456518 212 456524 264
rect 456576 252 456582 264
rect 467484 252 467512 552
rect 468846 484 468852 536
rect 468904 524 468910 536
rect 480714 524 480720 536
rect 468904 496 480720 524
rect 468904 484 468910 496
rect 480714 484 480720 496
rect 480772 484 480778 536
rect 485406 484 485412 536
rect 485464 524 485470 536
rect 498378 524 498384 536
rect 485464 496 498384 524
rect 485464 484 485470 496
rect 498378 484 498384 496
rect 498436 484 498442 536
rect 502794 484 502800 536
rect 502852 524 502858 536
rect 506032 524 506060 564
rect 517146 552 517152 564
rect 517204 552 517210 604
rect 518434 552 518440 604
rect 518492 552 518498 604
rect 518866 592 518894 632
rect 519446 620 519452 672
rect 519504 660 519510 672
rect 534810 660 534816 672
rect 519504 632 534816 660
rect 519504 620 519510 632
rect 534810 620 534816 632
rect 534868 620 534874 672
rect 529014 592 529020 604
rect 518866 564 529020 592
rect 529014 552 529020 564
rect 529072 552 529078 604
rect 533706 552 533712 604
rect 533764 552 533770 604
rect 534994 552 535000 604
rect 535052 552 535058 604
rect 535472 592 535500 700
rect 546678 688 546684 700
rect 546736 688 546742 740
rect 547846 700 551324 728
rect 536006 620 536012 672
rect 536064 660 536070 672
rect 547846 660 547874 700
rect 551186 660 551192 672
rect 536064 632 547874 660
rect 549916 632 551192 660
rect 536064 620 536070 632
rect 549070 592 549076 604
rect 535472 564 549076 592
rect 549070 552 549076 564
rect 549128 552 549134 604
rect 502852 496 506060 524
rect 502852 484 502858 496
rect 506106 484 506112 536
rect 506164 524 506170 536
rect 515766 524 515772 536
rect 506164 496 515772 524
rect 506164 484 506170 496
rect 515766 484 515772 496
rect 515824 484 515830 536
rect 518452 524 518480 552
rect 533724 524 533752 552
rect 518452 496 533752 524
rect 535012 524 535040 552
rect 549916 524 549944 632
rect 551186 620 551192 632
rect 551244 620 551250 672
rect 550266 552 550272 604
rect 550324 552 550330 604
rect 550358 552 550364 604
rect 550416 552 550422 604
rect 551296 592 551324 700
rect 551370 688 551376 740
rect 551428 728 551434 740
rect 569126 728 569132 740
rect 551428 700 569132 728
rect 551428 688 551434 700
rect 569126 688 569132 700
rect 569184 688 569190 740
rect 558086 620 558092 672
rect 558144 660 558150 672
rect 576302 660 576308 672
rect 558144 632 576308 660
rect 558144 620 558150 632
rect 576302 620 576308 632
rect 576360 620 576366 672
rect 552658 592 552664 604
rect 551296 564 552664 592
rect 552658 552 552664 564
rect 552716 552 552722 604
rect 568022 592 568028 604
rect 553964 564 568028 592
rect 535012 496 549944 524
rect 479702 416 479708 468
rect 479760 456 479766 468
rect 492490 456 492496 468
rect 479760 428 492496 456
rect 479760 416 479766 428
rect 492490 416 492496 428
rect 492548 416 492554 468
rect 496262 416 496268 468
rect 496320 456 496326 468
rect 509878 456 509884 468
rect 496320 428 509884 456
rect 496320 416 496326 428
rect 509878 416 509884 428
rect 509936 416 509942 468
rect 512822 416 512828 468
rect 512880 456 512886 468
rect 528002 456 528008 468
rect 512880 428 528008 456
rect 512880 416 512886 428
rect 528002 416 528008 428
rect 528060 416 528066 468
rect 529382 416 529388 468
rect 529440 456 529446 468
rect 545666 456 545672 468
rect 529440 428 545672 456
rect 529440 416 529446 428
rect 545666 416 545672 428
rect 545724 416 545730 468
rect 550284 456 550312 552
rect 550376 524 550404 552
rect 553964 524 553992 564
rect 568022 552 568028 564
rect 568080 552 568086 604
rect 575106 552 575112 604
rect 575164 552 575170 604
rect 550376 496 553992 524
rect 556982 484 556988 536
rect 557040 524 557046 536
rect 575124 524 575152 552
rect 557040 496 575152 524
rect 557040 484 557046 496
rect 567010 456 567016 468
rect 547846 428 550312 456
rect 553412 428 567016 456
rect 467650 348 467656 400
rect 467708 388 467714 400
rect 479150 388 479156 400
rect 467708 360 479156 388
rect 467708 348 467714 360
rect 479150 348 479156 360
rect 479208 348 479214 400
rect 484210 348 484216 400
rect 484268 388 484274 400
rect 497274 388 497280 400
rect 484268 360 497280 388
rect 484268 348 484274 360
rect 497274 348 497280 360
rect 497332 348 497338 400
rect 500770 348 500776 400
rect 500828 388 500834 400
rect 514938 388 514944 400
rect 500828 360 514944 388
rect 500828 348 500834 360
rect 514938 348 514944 360
rect 514996 348 515002 400
rect 516134 348 516140 400
rect 516192 388 516198 400
rect 531498 388 531504 400
rect 516192 360 531504 388
rect 516192 348 516198 360
rect 531498 348 531504 360
rect 531556 348 531562 400
rect 533890 348 533896 400
rect 533948 388 533954 400
rect 547846 388 547874 428
rect 533948 360 547874 388
rect 533948 348 533954 360
rect 549254 348 549260 400
rect 549312 388 549318 400
rect 553412 388 553440 428
rect 567010 416 567016 428
rect 567068 416 567074 468
rect 549312 360 553440 388
rect 549312 348 549318 360
rect 555878 348 555884 400
rect 555936 388 555942 400
rect 573726 388 573732 400
rect 555936 360 573732 388
rect 555936 348 555942 360
rect 573726 348 573732 360
rect 573784 348 573790 400
rect 473078 280 473084 332
rect 473136 320 473142 332
rect 485038 320 485044 332
rect 473136 292 485044 320
rect 473136 280 473142 292
rect 485038 280 485044 292
rect 485096 280 485102 332
rect 485498 280 485504 332
rect 485556 320 485562 332
rect 495710 320 495716 332
rect 485556 292 495716 320
rect 485556 280 485562 292
rect 495710 280 495716 292
rect 495768 280 495774 332
rect 499574 280 499580 332
rect 499632 320 499638 332
rect 513374 320 513380 332
rect 499632 292 513380 320
rect 499632 280 499638 292
rect 513374 280 513380 292
rect 513432 280 513438 332
rect 522758 280 522764 332
rect 522816 320 522822 332
rect 538214 320 538220 332
rect 522816 292 538220 320
rect 522816 280 522822 292
rect 538214 280 538220 292
rect 538272 280 538278 332
rect 539318 280 539324 332
rect 539376 320 539382 332
rect 556338 320 556344 332
rect 539376 292 556344 320
rect 539376 280 539382 292
rect 556338 280 556344 292
rect 556396 280 556402 332
rect 556430 280 556436 332
rect 556488 320 556494 332
rect 558730 320 558736 332
rect 556488 292 558736 320
rect 556488 280 556494 292
rect 558730 280 558736 292
rect 558788 280 558794 332
rect 560202 280 560208 332
rect 560260 320 560266 332
rect 578786 320 578792 332
rect 560260 292 578792 320
rect 560260 280 560266 292
rect 578786 280 578792 292
rect 578844 280 578850 332
rect 456576 224 467512 252
rect 456576 212 456582 224
rect 471882 212 471888 264
rect 471940 252 471946 264
rect 483842 252 483848 264
rect 471940 224 483848 252
rect 471940 212 471946 224
rect 483842 212 483848 224
rect 483900 212 483906 264
rect 488442 212 488448 264
rect 488500 252 488506 264
rect 501598 252 501604 264
rect 488500 224 501604 252
rect 488500 212 488506 224
rect 501598 212 501604 224
rect 501656 212 501662 264
rect 505002 212 505008 264
rect 505060 252 505066 264
rect 519722 252 519728 264
rect 505060 224 519728 252
rect 505060 212 505066 224
rect 519722 212 519728 224
rect 519780 212 519786 264
rect 521562 212 521568 264
rect 521620 252 521626 264
rect 537386 252 537392 264
rect 521620 224 537392 252
rect 521620 212 521626 224
rect 537386 212 537392 224
rect 537444 212 537450 264
rect 538122 212 538128 264
rect 538180 252 538186 264
rect 554774 252 554780 264
rect 538180 224 554780 252
rect 538180 212 538186 224
rect 554774 212 554780 224
rect 554832 212 554838 264
rect 563606 212 563612 264
rect 563664 252 563670 264
rect 583570 252 583576 264
rect 563664 224 583576 252
rect 563664 212 563670 224
rect 583570 212 583576 224
rect 583628 212 583634 264
rect 223482 184 223488 196
rect 218072 156 223488 184
rect 223482 144 223488 156
rect 223540 144 223546 196
rect 381446 144 381452 196
rect 381504 184 381510 196
rect 386966 184 386972 196
rect 381504 156 386972 184
rect 381504 144 381510 156
rect 386966 144 386972 156
rect 387024 144 387030 196
rect 399938 144 399944 196
rect 399996 184 400002 196
rect 407022 184 407028 196
rect 399996 156 407028 184
rect 399996 144 400002 156
rect 407022 144 407028 156
rect 407080 144 407086 196
rect 411162 144 411168 196
rect 411220 184 411226 196
rect 418798 184 418804 196
rect 411220 156 418804 184
rect 411220 144 411226 156
rect 418798 144 418804 156
rect 418856 144 418862 196
rect 422202 144 422208 196
rect 422260 184 422266 196
rect 431034 184 431040 196
rect 422260 156 431040 184
rect 422260 144 422266 156
rect 431034 144 431040 156
rect 431092 144 431098 196
rect 433058 144 433064 196
rect 433116 184 433122 196
rect 442810 184 442816 196
rect 433116 156 442816 184
rect 433116 144 433122 156
rect 442810 144 442816 156
rect 442868 144 442874 196
rect 444282 144 444288 196
rect 444340 184 444346 196
rect 454310 184 454316 196
rect 444340 156 454316 184
rect 444340 144 444346 156
rect 454310 144 454316 156
rect 454368 144 454374 196
rect 455322 144 455328 196
rect 455380 184 455386 196
rect 466086 184 466092 196
rect 455380 156 466092 184
rect 455380 144 455386 156
rect 466086 144 466092 156
rect 466144 144 466150 196
rect 466454 144 466460 196
rect 466512 184 466518 196
rect 478322 184 478328 196
rect 466512 156 478328 184
rect 466512 144 466518 156
rect 478322 144 478328 156
rect 478380 144 478386 196
rect 488626 144 488632 196
rect 488684 184 488690 196
rect 490926 184 490932 196
rect 488684 156 490932 184
rect 488684 144 488690 156
rect 490926 144 490932 156
rect 490984 144 490990 196
rect 495158 144 495164 196
rect 495216 184 495222 196
rect 509050 184 509056 196
rect 495216 156 509056 184
rect 495216 144 495222 156
rect 509050 144 509056 156
rect 509108 144 509114 196
rect 511718 144 511724 196
rect 511776 184 511782 196
rect 526438 184 526444 196
rect 511776 156 526444 184
rect 511776 144 511782 156
rect 526438 144 526444 156
rect 526496 144 526502 196
rect 528278 144 528284 196
rect 528336 184 528342 196
rect 544562 184 544568 196
rect 528336 156 544568 184
rect 528336 144 528342 156
rect 544562 144 544568 156
rect 544620 144 544626 196
rect 544838 144 544844 196
rect 544896 184 544902 196
rect 562226 184 562232 196
rect 544896 156 562232 184
rect 544896 144 544902 156
rect 562226 144 562232 156
rect 562284 144 562290 196
rect 562502 144 562508 196
rect 562560 184 562566 196
rect 582006 184 582012 196
rect 562560 156 582012 184
rect 562560 144 562566 156
rect 582006 144 582012 156
rect 582064 144 582070 196
rect 382 76 388 128
rect 440 116 446 128
rect 20346 116 20352 128
rect 440 88 20352 116
rect 440 76 446 88
rect 20346 76 20352 88
rect 20404 76 20410 128
rect 38010 116 38016 128
rect 26206 88 38016 116
rect 19610 8 19616 60
rect 19668 48 19674 60
rect 26206 48 26234 88
rect 38010 76 38016 88
rect 38068 76 38074 128
rect 38562 76 38568 128
rect 38620 116 38626 128
rect 55674 116 55680 128
rect 38620 88 55680 116
rect 38620 76 38626 88
rect 55674 76 55680 88
rect 55732 76 55738 128
rect 57054 76 57060 128
rect 57112 116 57118 128
rect 73338 116 73344 128
rect 57112 88 73344 116
rect 57112 76 57118 88
rect 73338 76 73344 88
rect 73396 76 73402 128
rect 75178 76 75184 128
rect 75236 116 75242 128
rect 89898 116 89904 128
rect 75236 88 89904 116
rect 75236 76 75242 88
rect 89898 76 89904 88
rect 89956 76 89962 128
rect 90174 76 90180 128
rect 90232 116 90238 128
rect 104250 116 104256 128
rect 90232 88 104256 116
rect 90232 76 90238 88
rect 104250 76 104256 88
rect 104308 76 104314 128
rect 104342 76 104348 128
rect 104400 116 104406 128
rect 117406 116 117412 128
rect 104400 88 117412 116
rect 104400 76 104406 88
rect 117406 76 117412 88
rect 117464 76 117470 128
rect 120902 76 120908 128
rect 120960 116 120966 128
rect 132770 116 132776 128
rect 120960 88 132776 116
rect 120960 76 120966 88
rect 132770 76 132776 88
rect 132828 76 132834 128
rect 134334 76 134340 128
rect 134392 116 134398 128
rect 145098 116 145104 128
rect 134392 88 145104 116
rect 134392 76 134398 88
rect 145098 76 145104 88
rect 145156 76 145162 128
rect 157242 116 157248 128
rect 147646 88 157248 116
rect 19668 20 26234 48
rect 19668 8 19674 20
rect 147306 8 147312 60
rect 147364 48 147370 60
rect 147646 48 147674 88
rect 157242 76 157248 88
rect 157300 76 157306 128
rect 157978 76 157984 128
rect 158036 116 158042 128
rect 167362 116 167368 128
rect 158036 88 167368 116
rect 158036 76 158042 88
rect 167362 76 167368 88
rect 167420 76 167426 128
rect 168650 76 168656 128
rect 168708 116 168714 128
rect 177114 116 177120 128
rect 168708 88 177120 116
rect 168708 76 168714 88
rect 177114 76 177120 88
rect 177172 76 177178 128
rect 180426 76 180432 128
rect 180484 116 180490 128
rect 188154 116 188160 128
rect 180484 88 188160 116
rect 180484 76 180490 88
rect 188154 76 188160 88
rect 188212 76 188218 128
rect 228542 76 228548 128
rect 228600 116 228606 128
rect 232498 116 232504 128
rect 228600 88 232504 116
rect 228600 76 228606 88
rect 232498 76 232504 88
rect 232556 76 232562 128
rect 344922 76 344928 128
rect 344980 116 344986 128
rect 348234 116 348240 128
rect 344980 88 348240 116
rect 344980 76 344986 88
rect 348234 76 348240 88
rect 348292 76 348298 128
rect 372522 76 372528 128
rect 372580 116 372586 128
rect 377858 116 377864 128
rect 372580 88 377864 116
rect 372580 76 372586 88
rect 377858 76 377864 88
rect 377916 76 377922 128
rect 383378 76 383384 128
rect 383436 116 383442 128
rect 389634 116 389640 128
rect 383436 88 389640 116
rect 383436 76 383442 88
rect 389634 76 389640 88
rect 389692 76 389698 128
rect 405642 76 405648 128
rect 405700 116 405706 128
rect 412910 116 412916 128
rect 405700 88 412916 116
rect 405700 76 405706 88
rect 412910 76 412916 88
rect 412968 76 412974 128
rect 413462 76 413468 128
rect 413520 116 413526 128
rect 421190 116 421196 128
rect 413520 88 421196 116
rect 413520 76 413526 88
rect 421190 76 421196 88
rect 421248 76 421254 128
rect 427722 76 427728 128
rect 427780 116 427786 128
rect 436922 116 436928 128
rect 427780 88 436928 116
rect 427780 76 427786 88
rect 436922 76 436928 88
rect 436980 76 436986 128
rect 438762 76 438768 128
rect 438820 116 438826 128
rect 448422 116 448428 128
rect 438820 88 448428 116
rect 438820 76 438826 88
rect 448422 76 448428 88
rect 448480 76 448486 128
rect 449618 76 449624 128
rect 449676 116 449682 128
rect 460198 116 460204 128
rect 449676 88 460204 116
rect 449676 76 449682 88
rect 460198 76 460204 88
rect 460256 76 460262 128
rect 460842 76 460848 128
rect 460900 116 460906 128
rect 472434 116 472440 128
rect 460900 88 472440 116
rect 460900 76 460906 88
rect 472434 76 472440 88
rect 472492 76 472498 128
rect 477402 76 477408 128
rect 477460 116 477466 128
rect 490098 116 490104 128
rect 477460 88 490104 116
rect 477460 76 477466 88
rect 490098 76 490104 88
rect 490156 76 490162 128
rect 493962 76 493968 128
rect 494020 116 494026 128
rect 507486 116 507492 128
rect 494020 88 507492 116
rect 494020 76 494026 88
rect 507486 76 507492 88
rect 507544 76 507550 128
rect 510522 76 510528 128
rect 510580 116 510586 128
rect 525610 116 525616 128
rect 510580 88 525616 116
rect 510580 76 510586 88
rect 525610 76 525616 88
rect 525668 76 525674 128
rect 527082 76 527088 128
rect 527140 116 527146 128
rect 542998 116 543004 128
rect 527140 88 543004 116
rect 527140 76 527146 88
rect 542998 76 543004 88
rect 543056 76 543062 128
rect 543642 76 543648 128
rect 543700 116 543706 128
rect 560662 116 560668 128
rect 543700 88 560668 116
rect 543700 76 543706 88
rect 560662 76 560668 88
rect 560720 76 560726 128
rect 561398 76 561404 128
rect 561456 116 561462 128
rect 581178 116 581184 128
rect 561456 88 581184 116
rect 561456 76 561462 88
rect 581178 76 581184 88
rect 581236 76 581242 128
rect 147364 20 147674 48
rect 147364 8 147370 20
rect 151998 8 152004 60
rect 152056 48 152062 60
rect 161658 48 161664 60
rect 152056 20 161664 48
rect 152056 8 152062 20
rect 161658 8 161664 20
rect 161716 8 161722 60
rect 467282 8 467288 60
rect 467340 48 467346 60
rect 470042 48 470048 60
rect 467340 20 470048 48
rect 467340 8 467346 20
rect 470042 8 470048 20
rect 470100 8 470106 60
<< via1 >>
rect 59176 2864 59228 2916
rect 64558 2864 64610 2916
rect 67640 2864 67692 2916
rect 70078 2864 70130 2916
rect 71780 2864 71832 2916
rect 74494 2864 74546 2916
rect 75460 2864 75512 2916
rect 76702 2864 76754 2916
rect 80152 2864 80204 2916
rect 84430 2864 84482 2916
rect 85396 2864 85448 2916
rect 86638 2864 86690 2916
rect 86776 2864 86828 2916
rect 87742 2864 87794 2916
rect 88156 2864 88208 2916
rect 92158 2864 92210 2916
rect 92480 2864 92532 2916
rect 94366 2864 94418 2916
rect 94596 2864 94648 2916
rect 95470 2864 95522 2916
rect 95700 2864 95752 2916
rect 97678 2864 97730 2916
rect 98000 2864 98052 2916
rect 100990 2864 101042 2916
rect 102232 2864 102284 2916
rect 105406 2864 105458 2916
rect 105544 2864 105596 2916
rect 106510 2864 106562 2916
rect 107752 2864 107804 2916
rect 109822 2864 109874 2916
rect 110420 2864 110472 2916
rect 113134 2864 113186 2916
rect 114744 2864 114796 2916
rect 116446 2864 116498 2916
rect 117320 2864 117372 2916
rect 119758 2864 119810 2916
rect 120080 2864 120132 2916
rect 124174 2864 124226 2916
rect 125140 2864 125192 2916
rect 127486 2864 127538 2916
rect 127624 2864 127676 2916
rect 129694 2864 129746 2916
rect 133236 2864 133288 2916
rect 134110 2864 134162 2916
rect 136640 2864 136692 2916
rect 139630 2864 139682 2916
rect 144184 2864 144236 2916
rect 146254 2864 146306 2916
rect 149060 2864 149112 2916
rect 151774 2864 151826 2916
rect 153384 2864 153436 2916
rect 155086 2864 155138 2916
rect 155960 2864 156012 2916
rect 158398 2864 158450 2916
rect 158720 2864 158772 2916
rect 162814 2864 162866 2916
rect 167000 2864 167052 2916
rect 169438 2864 169490 2916
rect 169576 2864 169628 2916
rect 170542 2864 170594 2916
rect 172980 2864 173032 2916
rect 174958 2864 175010 2916
rect 175280 2864 175332 2916
rect 178270 2864 178322 2916
rect 179512 2864 179564 2916
rect 181582 2864 181634 2916
rect 181720 2864 181772 2916
rect 182686 2864 182738 2916
rect 187700 2864 187752 2916
rect 189310 2864 189362 2916
rect 205640 2864 205692 2916
rect 208078 2864 208130 2916
rect 211620 2864 211672 2916
rect 213598 2864 213650 2916
rect 213736 2864 213788 2916
rect 214702 2864 214754 2916
rect 214840 2864 214892 2916
rect 215806 2864 215858 2916
rect 216680 2864 216732 2916
rect 219118 2864 219170 2916
rect 220360 2864 220412 2916
rect 221326 2864 221378 2916
rect 221464 2864 221516 2916
rect 222430 2864 222482 2916
rect 222568 2864 222620 2916
rect 224638 2864 224690 2916
rect 224776 2864 224828 2916
rect 225742 2864 225794 2916
rect 226524 2864 226576 2916
rect 227950 2864 228002 2916
rect 230572 2864 230624 2916
rect 232366 2864 232418 2916
rect 232504 2864 232556 2916
rect 233470 2864 233522 2916
rect 234712 2864 234764 2916
rect 236782 2864 236834 2916
rect 242900 2864 242952 2916
rect 246718 2864 246770 2916
rect 247592 2864 247644 2916
rect 251134 2864 251186 2916
rect 253480 2864 253532 2916
rect 256654 2864 256706 2916
rect 257068 2864 257120 2916
rect 259966 2864 260018 2916
rect 261760 2864 261812 2916
rect 264382 2864 264434 2916
rect 265348 2864 265400 2916
rect 267694 2864 267746 2916
rect 267832 2864 267884 2916
rect 269902 2864 269954 2916
rect 271236 2864 271288 2916
rect 273214 2864 273266 2916
rect 273628 2864 273680 2916
rect 275422 2864 275474 2916
rect 276020 2864 276072 2916
rect 277630 2864 277682 2916
rect 278320 2864 278372 2916
rect 279838 2864 279890 2916
rect 280712 2864 280764 2916
rect 282046 2864 282098 2916
rect 283150 2864 283202 2916
rect 286600 2864 286652 2916
rect 287566 2864 287618 2916
rect 287796 2864 287848 2916
rect 288670 2864 288722 2916
rect 293684 2864 293736 2916
rect 294190 2864 294242 2916
rect 320686 2864 320738 2916
rect 322112 2864 322164 2916
rect 322894 2864 322946 2916
rect 324412 2864 324464 2916
rect 325102 2864 325154 2916
rect 326804 2864 326856 2916
rect 329518 2864 329570 2916
rect 331588 2864 331640 2916
rect 331726 2864 331778 2916
rect 333796 2864 333848 2916
rect 335038 2864 335090 2916
rect 336464 2864 336516 2916
rect 340558 2864 340610 2916
rect 343364 2864 343416 2916
rect 346078 2864 346130 2916
rect 347596 2864 347648 2916
rect 348286 2864 348338 2916
rect 349896 2864 349948 2916
rect 352702 2864 352754 2916
rect 355784 2864 355836 2916
rect 358222 2864 358274 2916
rect 360108 2864 360160 2916
rect 362638 2864 362690 2916
rect 363512 2864 363564 2916
rect 363742 2864 363794 2916
rect 366180 2864 366232 2916
rect 369262 2864 369314 2916
rect 370228 2864 370280 2916
rect 370366 2864 370418 2916
rect 372712 2864 372764 2916
rect 373678 2864 373730 2916
rect 375104 2864 375156 2916
rect 375886 2864 375938 2916
rect 378508 2864 378560 2916
rect 379198 2864 379250 2916
rect 380164 2864 380216 2916
rect 380302 2864 380354 2916
rect 382280 2864 382332 2916
rect 386926 2864 386978 2916
rect 387892 2864 387944 2916
rect 388030 2864 388082 2916
rect 390652 2864 390704 2916
rect 391342 2864 391394 2916
rect 394424 2864 394476 2916
rect 396862 2864 396914 2916
rect 398748 2864 398800 2916
rect 399070 2864 399122 2916
rect 401600 2864 401652 2916
rect 402382 2864 402434 2916
rect 404268 2864 404320 2916
rect 406798 2864 406850 2916
rect 407764 2864 407816 2916
rect 407902 2864 407954 2916
rect 409788 2864 409840 2916
rect 415630 2864 415682 2916
rect 423772 2864 423824 2916
rect 424462 2864 424514 2916
rect 425428 2864 425480 2916
rect 425566 2864 425618 2916
rect 428740 2864 428792 2916
rect 428878 2864 428930 2916
rect 429844 2864 429896 2916
rect 429982 2864 430034 2916
rect 433156 2864 433208 2916
rect 439918 2864 439970 2916
rect 442908 2864 442960 2916
rect 450958 2864 451010 2916
rect 452568 2864 452620 2916
rect 461998 2864 462050 2916
rect 63500 2796 63552 2848
rect 67870 2796 67922 2848
rect 73160 2796 73212 2848
rect 75598 2796 75650 2848
rect 76840 2796 76892 2848
rect 81118 2796 81170 2848
rect 100760 2796 100812 2848
rect 103198 2796 103250 2848
rect 150440 2796 150492 2848
rect 152878 2796 152930 2848
rect 204260 2796 204312 2848
rect 206974 2796 207026 2848
rect 215300 2796 215352 2848
rect 217968 2796 218020 2848
rect 218060 2796 218112 2848
rect 220222 2796 220274 2848
rect 224960 2796 225012 2848
rect 226846 2796 226898 2848
rect 249892 2796 249944 2848
rect 253342 2796 253394 2848
rect 259460 2796 259512 2848
rect 262174 2796 262226 2848
rect 266544 2796 266596 2848
rect 268798 2796 268850 2848
rect 272432 2796 272484 2848
rect 274318 2796 274370 2848
rect 274824 2796 274876 2848
rect 276526 2796 276578 2848
rect 279516 2796 279568 2848
rect 280942 2796 280994 2848
rect 281908 2796 281960 2848
rect 285404 2796 285456 2848
rect 286462 2796 286514 2848
rect 316270 2796 316322 2848
rect 317328 2796 317380 2848
rect 336142 2796 336194 2848
rect 338672 2796 338724 2848
rect 342766 2796 342818 2848
rect 345756 2796 345808 2848
rect 347182 2796 347234 2848
rect 348792 2796 348844 2848
rect 349390 2796 349442 2848
rect 352840 2796 352892 2848
rect 354910 2796 354962 2848
rect 358728 2796 358780 2848
rect 359326 2796 359378 2848
rect 362500 2796 362552 2848
rect 365950 2796 366002 2848
rect 369768 2796 369820 2848
rect 374782 2796 374834 2848
rect 376668 2796 376720 2848
rect 382510 2796 382562 2848
rect 387708 2796 387760 2848
rect 393550 2796 393602 2848
rect 396724 2796 396776 2848
rect 397966 2796 398018 2848
rect 399852 2796 399904 2848
rect 403486 2796 403538 2848
rect 407028 2796 407080 2848
rect 409006 2796 409058 2848
rect 416596 2796 416648 2848
rect 432190 2796 432242 2848
rect 438952 2796 439004 2848
rect 442126 2796 442178 2848
rect 451188 2796 451240 2848
rect 452062 2796 452114 2848
rect 462228 2796 462280 2848
rect 463102 2864 463154 2916
rect 464068 2864 464120 2916
rect 464206 2864 464258 2916
rect 466184 2864 466236 2916
rect 476350 2864 476402 2916
rect 478328 2864 478380 2916
rect 490702 2864 490754 2916
rect 492588 2864 492640 2916
rect 506158 2864 506210 2916
rect 507860 2864 507912 2916
rect 508366 2864 508418 2916
rect 509976 2864 510028 2916
rect 523822 2864 523874 2916
rect 525708 2864 525760 2916
rect 540382 2864 540434 2916
rect 541348 2864 541400 2916
rect 541486 2864 541538 2916
rect 556436 2864 556488 2916
rect 463608 2796 463660 2848
rect 465310 2796 465362 2848
rect 476948 2796 477000 2848
rect 478558 2796 478610 2848
rect 488632 2796 488684 2848
rect 491806 2796 491858 2848
rect 505376 2796 505428 2848
rect 509470 2796 509522 2848
rect 524236 2796 524288 2848
rect 524926 2796 524978 2848
rect 540796 2796 540848 2848
rect 28908 1300 28960 1352
rect 23020 1232 23072 1284
rect 17040 1096 17092 1148
rect 18236 1028 18288 1080
rect 35992 1232 36044 1284
rect 53472 1232 53524 1284
rect 31484 1164 31536 1216
rect 44640 1164 44692 1216
rect 51356 1164 51408 1216
rect 46848 1096 46900 1148
rect 18880 960 18932 1012
rect 22560 960 22612 1012
rect 41328 1028 41380 1080
rect 46664 1028 46716 1080
rect 21180 892 21232 944
rect 25872 892 25924 944
rect 35808 960 35860 1012
rect 40684 960 40736 1012
rect 36912 892 36964 944
rect 47216 960 47268 1012
rect 54576 960 54628 1012
rect 65524 1164 65576 1216
rect 58440 1096 58492 1148
rect 71780 1096 71832 1148
rect 76840 1096 76892 1148
rect 77392 1096 77444 1148
rect 88156 1096 88208 1148
rect 63500 1028 63552 1080
rect 69112 1028 69164 1080
rect 80152 1028 80204 1080
rect 97448 1028 97500 1080
rect 110880 1028 110932 1080
rect 63408 960 63460 1012
rect 71504 960 71556 1012
rect 85396 960 85448 1012
rect 91560 960 91612 1012
rect 102232 960 102284 1012
rect 57888 892 57940 944
rect 59636 892 59688 944
rect 73160 892 73212 944
rect 83280 892 83332 944
rect 11152 824 11204 876
rect 30288 824 30340 876
rect 30380 824 30432 876
rect 47952 824 48004 876
rect 12348 756 12400 808
rect 31392 756 31444 808
rect 34796 756 34848 808
rect 52368 756 52420 808
rect 13544 688 13596 740
rect 32496 688 32548 740
rect 41880 688 41932 740
rect 5264 620 5316 672
rect 24768 620 24820 672
rect 6460 552 6512 604
rect 21180 552 21232 604
rect 24216 552 24268 604
rect 42432 620 42484 672
rect 25320 552 25372 604
rect 43536 620 43588 672
rect 47860 688 47912 740
rect 59176 824 59228 876
rect 60832 824 60884 876
rect 53748 756 53800 808
rect 67640 756 67692 808
rect 52552 688 52604 740
rect 68928 688 68980 740
rect 58992 620 59044 672
rect 64328 620 64380 672
rect 76932 824 76984 876
rect 82176 824 82228 876
rect 86868 892 86920 944
rect 98000 892 98052 944
rect 95700 824 95752 876
rect 100760 892 100812 944
rect 105728 892 105780 944
rect 118608 1164 118660 1216
rect 537116 1164 537168 1216
rect 553768 1164 553820 1216
rect 72608 756 72660 808
rect 86776 756 86828 808
rect 89168 756 89220 808
rect 99840 824 99892 876
rect 110420 824 110472 876
rect 70308 688 70360 740
rect 85488 688 85540 740
rect 87972 688 88024 740
rect 102048 756 102100 808
rect 106004 756 106056 808
rect 107752 756 107804 808
rect 96252 688 96304 740
rect 43076 552 43128 604
rect 60096 552 60148 604
rect 62028 552 62080 604
rect 75460 620 75512 672
rect 76196 620 76248 672
rect 91008 620 91060 672
rect 95148 620 95200 672
rect 14556 484 14608 536
rect 33416 484 33468 536
rect 37004 484 37056 536
rect 47216 484 47268 536
rect 7840 416 7892 468
rect 26976 416 27028 468
rect 31116 416 31168 468
rect 49148 484 49200 536
rect 77760 484 77812 536
rect 48780 416 48832 468
rect 65708 416 65760 468
rect 66904 416 66956 468
rect 76932 416 76984 468
rect 79692 552 79744 604
rect 82084 552 82136 604
rect 96528 552 96580 604
rect 101036 552 101088 604
rect 92480 484 92532 536
rect 79968 416 80020 468
rect 84660 416 84712 468
rect 98828 416 98880 468
rect 103336 688 103388 740
rect 114744 1096 114796 1148
rect 541348 1096 541400 1148
rect 557356 1096 557408 1148
rect 111616 1028 111668 1080
rect 101312 620 101364 672
rect 107568 620 107620 672
rect 117320 892 117372 944
rect 509976 1028 510028 1080
rect 523040 1028 523092 1080
rect 525708 1028 525760 1080
rect 539600 1028 539652 1080
rect 548156 1028 548208 1080
rect 565636 1028 565688 1080
rect 143448 960 143500 1012
rect 149060 960 149112 1012
rect 470876 960 470928 1012
rect 482836 960 482888 1012
rect 487436 960 487488 1012
rect 500592 960 500644 1012
rect 501788 960 501840 1012
rect 506112 960 506164 1012
rect 507860 960 507912 1012
rect 120080 892 120132 944
rect 127532 892 127584 944
rect 133236 892 133288 944
rect 135260 892 135312 944
rect 144184 892 144236 944
rect 148324 892 148376 944
rect 155960 892 156012 944
rect 190828 892 190880 944
rect 198096 892 198148 944
rect 466184 892 466236 944
rect 475752 892 475804 944
rect 478328 892 478380 944
rect 488816 892 488868 944
rect 492588 892 492640 944
rect 115204 824 115256 876
rect 125140 824 125192 876
rect 128176 824 128228 876
rect 136640 824 136692 876
rect 140044 824 140096 876
rect 150624 824 150676 876
rect 161480 824 161532 876
rect 169576 824 169628 876
rect 183744 824 183796 876
rect 191472 824 191524 876
rect 210976 824 211028 876
rect 216864 824 216916 876
rect 433064 824 433116 876
rect 433248 824 433300 876
rect 464068 824 464120 876
rect 474556 824 474608 876
rect 475292 824 475344 876
rect 487620 824 487672 876
rect 492956 824 493008 876
rect 503996 892 504048 944
rect 518256 892 518308 944
rect 520556 960 520608 1012
rect 536104 960 536156 1012
rect 547052 960 547104 1012
rect 564440 960 564492 1012
rect 520740 892 520792 944
rect 526076 892 526128 944
rect 541992 892 542044 944
rect 545948 892 546000 944
rect 563244 892 563296 944
rect 112812 756 112864 808
rect 106004 552 106056 604
rect 8944 348 8996 400
rect 9772 280 9824 332
rect 21180 280 21232 332
rect 1492 212 1544 264
rect 21364 348 21416 400
rect 26332 348 26384 400
rect 31484 348 31536 400
rect 32220 348 32272 400
rect 49976 348 50028 400
rect 55128 348 55180 400
rect 71136 348 71188 400
rect 78404 348 78456 400
rect 29184 280 29236 332
rect 33784 280 33836 332
rect 51172 280 51224 332
rect 56232 280 56284 332
rect 72240 280 72292 332
rect 73620 280 73672 332
rect 88800 280 88852 332
rect 92572 348 92624 400
rect 105544 348 105596 400
rect 93216 280 93268 332
rect 94136 280 94188 332
rect 101312 280 101364 332
rect 106740 484 106792 536
rect 108120 552 108172 604
rect 108672 348 108724 400
rect 114192 484 114244 536
rect 123484 756 123536 808
rect 117596 688 117648 740
rect 127624 688 127676 740
rect 129372 756 129424 808
rect 140688 756 140740 808
rect 141240 756 141292 808
rect 143448 756 143500 808
rect 143540 756 143592 808
rect 153936 756 153988 808
rect 164884 756 164936 808
rect 173808 756 173860 808
rect 184940 756 184992 808
rect 192576 756 192628 808
rect 193220 756 193272 808
rect 200304 756 200356 808
rect 203892 756 203944 808
rect 210240 756 210292 808
rect 214472 756 214524 808
rect 218060 756 218112 808
rect 223948 756 224000 808
rect 229008 756 229060 808
rect 229836 756 229888 808
rect 234528 756 234580 808
rect 351644 756 351696 808
rect 355232 756 355284 808
rect 367008 756 367060 808
rect 371700 756 371752 808
rect 378048 756 378100 808
rect 383568 756 383620 808
rect 385868 756 385920 808
rect 391848 756 391900 808
rect 394516 756 394568 808
rect 401324 756 401376 808
rect 404636 756 404688 808
rect 411904 756 411956 808
rect 416688 756 416740 808
rect 424968 756 425020 808
rect 433156 756 433208 808
rect 439136 756 439188 808
rect 443276 756 443328 808
rect 451096 756 451148 808
rect 135168 688 135220 740
rect 144736 688 144788 740
rect 153384 688 153436 740
rect 166172 688 166224 740
rect 172980 688 173032 740
rect 173164 688 173216 740
rect 179512 688 179564 740
rect 181444 688 181496 740
rect 187700 688 187752 740
rect 118792 620 118844 672
rect 130752 620 130804 672
rect 136456 620 136508 672
rect 147312 620 147364 672
rect 149520 620 149572 672
rect 159456 620 159508 672
rect 160100 620 160152 672
rect 167000 620 167052 672
rect 167184 620 167236 672
rect 125232 552 125284 604
rect 130568 552 130620 604
rect 141792 552 141844 604
rect 142436 552 142488 604
rect 150440 552 150492 604
rect 150624 552 150676 604
rect 154212 552 154264 604
rect 163872 552 163924 604
rect 120816 484 120868 536
rect 124864 484 124916 536
rect 136272 484 136324 536
rect 120080 416 120132 468
rect 109132 348 109184 400
rect 121920 348 121972 400
rect 122472 348 122524 400
rect 127532 348 127584 400
rect 131580 416 131632 468
rect 142896 416 142948 468
rect 145748 416 145800 468
rect 131948 348 132000 400
rect 137468 348 137520 400
rect 148508 348 148560 400
rect 110696 280 110748 332
rect 123024 280 123076 332
rect 125692 280 125744 332
rect 137376 280 137428 332
rect 139032 280 139084 332
rect 149336 280 149388 332
rect 3056 144 3108 196
rect 18880 144 18932 196
rect 28080 212 28132 264
rect 44456 212 44508 264
rect 61200 212 61252 264
rect 63408 212 63460 264
rect 78864 212 78916 264
rect 81072 212 81124 264
rect 94596 212 94648 264
rect 98460 212 98512 264
rect 111984 212 112036 264
rect 114192 212 114244 264
rect 126336 212 126388 264
rect 126796 212 126848 264
rect 138480 212 138532 264
rect 21456 144 21508 196
rect 27896 144 27948 196
rect 45744 144 45796 196
rect 50344 144 50396 196
rect 66536 144 66588 196
rect 68192 144 68244 196
rect 83096 144 83148 196
rect 85856 144 85908 196
rect 99656 144 99708 196
rect 102416 144 102468 196
rect 115388 144 115440 196
rect 116584 144 116636 196
rect 128544 144 128596 196
rect 133144 144 133196 196
rect 144000 144 144052 196
rect 156420 416 156472 468
rect 165896 416 165948 468
rect 155592 348 155644 400
rect 165068 348 165120 400
rect 153200 280 153252 332
rect 158720 280 158772 332
rect 159088 280 159140 332
rect 168196 280 168248 332
rect 169576 620 169628 672
rect 175280 620 175332 672
rect 174268 552 174320 604
rect 181720 620 181772 672
rect 182548 620 182600 672
rect 190368 688 190420 740
rect 194416 688 194468 740
rect 201408 688 201460 740
rect 201500 688 201552 740
rect 205640 688 205692 740
rect 209780 688 209832 740
rect 214840 688 214892 740
rect 215668 688 215720 740
rect 220360 688 220412 740
rect 220452 688 220504 740
rect 224776 688 224828 740
rect 233424 688 233476 740
rect 237840 688 237892 740
rect 248788 688 248840 740
rect 252192 688 252244 740
rect 318524 688 318576 740
rect 319720 688 319772 740
rect 341708 688 341760 740
rect 344560 688 344612 740
rect 350448 688 350500 740
rect 354036 688 354088 740
rect 364892 688 364944 740
rect 369400 688 369452 740
rect 380164 688 380216 740
rect 384764 688 384816 740
rect 390652 688 390704 740
rect 394240 688 394292 740
rect 396724 688 396776 740
rect 400128 688 400180 740
rect 407764 688 407816 740
rect 414296 688 414348 740
rect 414572 688 414624 740
rect 422576 688 422628 740
rect 425428 688 425480 740
rect 433248 688 433300 740
rect 448796 688 448848 740
rect 459192 688 459244 740
rect 459836 688 459888 740
rect 471060 756 471112 808
rect 481916 756 481968 808
rect 494704 756 494756 808
rect 498476 756 498528 808
rect 503628 756 503680 808
rect 463608 688 463660 740
rect 188528 620 188580 672
rect 176660 552 176712 604
rect 184848 552 184900 604
rect 189724 552 189776 604
rect 195612 620 195664 672
rect 202512 620 202564 672
rect 195888 552 195940 604
rect 200304 552 200356 604
rect 204260 620 204312 672
rect 207388 620 207440 672
rect 211620 620 211672 672
rect 212172 620 212224 672
rect 215300 620 215352 672
rect 216864 620 216916 672
rect 221464 620 221516 672
rect 226340 620 226392 672
rect 231216 620 231268 672
rect 234620 620 234672 672
rect 238944 620 238996 672
rect 240508 620 240560 672
rect 244464 620 244516 672
rect 245200 620 245252 672
rect 248880 620 248932 672
rect 262956 620 263008 672
rect 265440 620 265492 672
rect 333980 620 334032 672
rect 336280 620 336332 672
rect 339500 620 339552 672
rect 342168 620 342220 672
rect 349896 620 349948 672
rect 351644 620 351696 672
rect 360476 620 360528 672
rect 364616 620 364668 672
rect 366180 620 366232 672
rect 368204 620 368256 672
rect 368296 620 368348 672
rect 372896 620 372948 672
rect 378508 620 378560 672
rect 381176 620 381228 672
rect 384672 620 384724 672
rect 202696 552 202748 604
rect 209136 552 209188 604
rect 213368 552 213420 604
rect 216680 552 216732 604
rect 218060 552 218112 604
rect 221556 552 221608 604
rect 224960 552 225012 604
rect 227536 552 227588 604
rect 230572 552 230624 604
rect 232228 552 232280 604
rect 234712 552 234764 604
rect 237012 552 237064 604
rect 241152 552 241204 604
rect 241704 552 241756 604
rect 245568 552 245620 604
rect 246396 552 246448 604
rect 250076 552 250128 604
rect 251180 552 251232 604
rect 254400 552 254452 604
rect 254676 552 254728 604
rect 257712 552 257764 604
rect 258264 552 258316 604
rect 261024 552 261076 604
rect 264152 552 264204 604
rect 266636 552 266688 604
rect 268844 552 268896 604
rect 270960 552 271012 604
rect 277124 552 277176 604
rect 278688 552 278740 604
rect 307484 552 307536 604
rect 307944 552 307996 604
rect 313004 552 313056 604
rect 313832 552 313884 604
rect 315212 552 315264 604
rect 316224 552 316276 604
rect 317236 552 317288 604
rect 318524 552 318576 604
rect 319628 552 319680 604
rect 320916 552 320968 604
rect 324044 552 324096 604
rect 325608 552 325660 604
rect 326252 552 326304 604
rect 328000 552 328052 604
rect 328368 552 328420 604
rect 330392 552 330444 604
rect 332876 552 332928 604
rect 335084 552 335136 604
rect 337292 552 337344 604
rect 339868 552 339920 604
rect 343916 552 343968 604
rect 346952 552 347004 604
rect 348792 552 348844 604
rect 350448 552 350500 604
rect 355784 552 355836 604
rect 356336 552 356388 604
rect 357164 552 357216 604
rect 361120 552 361172 604
rect 363512 552 363564 604
rect 367008 552 367060 604
rect 369768 552 369820 604
rect 370596 552 370648 604
rect 372712 552 372764 604
rect 375288 552 375340 604
rect 376668 552 376720 604
rect 379980 552 380032 604
rect 382280 552 382332 604
rect 385960 552 386012 604
rect 389088 620 389140 672
rect 395344 620 395396 672
rect 395804 620 395856 672
rect 390652 552 390704 604
rect 394424 552 394476 604
rect 397736 552 397788 604
rect 398748 620 398800 672
rect 403624 620 403676 672
rect 407028 620 407080 672
rect 410800 620 410852 672
rect 417792 620 417844 672
rect 402520 552 402572 604
rect 406016 552 406068 604
rect 409788 552 409840 604
rect 415492 552 415544 604
rect 417884 552 417936 604
rect 178040 484 178092 536
rect 185952 484 186004 536
rect 196992 484 197044 536
rect 172152 416 172204 468
rect 180432 416 180484 468
rect 192208 416 192260 468
rect 199292 416 199344 468
rect 170588 348 170640 400
rect 179328 348 179380 400
rect 196992 348 197044 400
rect 203616 348 203668 400
rect 208768 348 208820 400
rect 213736 348 213788 400
rect 176016 280 176068 332
rect 178868 280 178920 332
rect 187056 280 187108 332
rect 205272 280 205324 332
rect 211344 280 211396 332
rect 160560 212 160612 264
rect 162308 212 162360 264
rect 171600 212 171652 264
rect 186320 212 186372 264
rect 193680 212 193732 264
rect 198096 212 198148 264
rect 204720 212 204772 264
rect 206376 212 206428 264
rect 212448 212 212500 264
rect 156144 144 156196 196
rect 163872 144 163924 196
rect 172704 144 172756 196
rect 175648 144 175700 196
rect 183560 144 183612 196
rect 187148 144 187200 196
rect 194784 144 194836 196
rect 198924 144 198976 196
rect 205824 144 205876 196
rect 401600 484 401652 536
rect 225328 416 225380 468
rect 230112 416 230164 468
rect 239496 416 239548 468
rect 243360 416 243412 468
rect 361488 416 361540 468
rect 365628 416 365680 468
rect 371516 416 371568 468
rect 376300 416 376352 468
rect 377036 416 377088 468
rect 382188 416 382240 468
rect 387892 416 387944 468
rect 392860 416 392912 468
rect 219440 348 219492 400
rect 222568 348 222620 400
rect 222936 348 222988 400
rect 226524 348 226576 400
rect 231216 348 231268 400
rect 235632 348 235684 400
rect 236000 348 236052 400
rect 240048 348 240100 400
rect 244280 348 244332 400
rect 247776 348 247828 400
rect 252560 348 252612 400
rect 255504 348 255556 400
rect 256056 348 256108 400
rect 258816 348 258868 400
rect 260840 348 260892 400
rect 263232 348 263284 400
rect 270224 348 270276 400
rect 272064 348 272116 400
rect 311808 348 311860 400
rect 312452 348 312504 400
rect 314108 348 314160 400
rect 314844 348 314896 400
rect 321836 348 321888 400
rect 323124 348 323176 400
rect 327356 348 327408 400
rect 329012 348 329064 400
rect 330668 348 330720 400
rect 332508 348 332560 400
rect 336464 348 336516 400
rect 337292 348 337344 400
rect 338396 348 338448 400
rect 340788 348 340840 400
rect 347596 348 347648 400
rect 349068 348 349120 400
rect 355876 348 355928 400
rect 359740 348 359792 400
rect 360108 348 360160 400
rect 362132 348 362184 400
rect 362500 348 362552 400
rect 363696 348 363748 400
rect 370228 348 370280 400
rect 373908 348 373960 400
rect 375104 348 375156 400
rect 378692 348 378744 400
rect 392492 348 392544 400
rect 398748 348 398800 400
rect 399852 348 399904 400
rect 404636 348 404688 400
rect 404268 280 404320 332
rect 409420 280 409472 332
rect 410156 280 410208 332
rect 428740 620 428792 672
rect 434444 620 434496 672
rect 421196 552 421248 604
rect 429660 552 429712 604
rect 437940 620 437992 672
rect 438952 620 439004 672
rect 441528 620 441580 672
rect 442908 620 442960 672
rect 420000 416 420052 468
rect 428648 416 428700 468
rect 429844 416 429896 468
rect 435548 552 435600 604
rect 437756 552 437808 604
rect 447416 552 447468 604
rect 447692 620 447744 672
rect 458088 620 458140 672
rect 458732 620 458784 672
rect 467288 620 467340 672
rect 449808 552 449860 604
rect 450912 552 450964 604
rect 451188 552 451240 604
rect 452108 552 452160 604
rect 452568 552 452620 604
rect 461584 552 461636 604
rect 419172 348 419224 400
rect 427084 348 427136 400
rect 436560 484 436612 536
rect 446036 484 446088 536
rect 454316 484 454368 536
rect 464988 484 465040 536
rect 425980 280 426032 332
rect 426716 280 426768 332
rect 435732 348 435784 400
rect 445208 348 445260 400
rect 431132 280 431184 332
rect 440148 280 440200 332
rect 441068 280 441120 332
rect 451096 416 451148 468
rect 453488 416 453540 468
rect 457628 416 457680 468
rect 468576 620 468628 672
rect 467472 552 467524 604
rect 480812 688 480864 740
rect 493508 688 493560 740
rect 469772 620 469824 672
rect 481732 620 481784 672
rect 482928 620 482980 672
rect 485504 620 485556 672
rect 473452 552 473504 604
rect 474188 552 474240 604
rect 486332 620 486384 672
rect 499396 688 499448 740
rect 504180 824 504232 876
rect 507308 824 507360 876
rect 521844 824 521896 876
rect 531596 824 531648 876
rect 547880 824 547932 876
rect 552572 824 552624 876
rect 570328 824 570380 876
rect 503904 756 503956 808
rect 512460 756 512512 808
rect 517244 756 517296 808
rect 532332 756 532384 808
rect 506480 688 506532 740
rect 515036 688 515088 740
rect 530124 688 530176 740
rect 530492 688 530544 740
rect 532608 688 532660 740
rect 542636 756 542688 808
rect 559104 756 559156 808
rect 559196 756 559248 808
rect 577412 756 577464 808
rect 497372 620 497424 672
rect 511264 620 511316 672
rect 513932 620 513984 672
rect 486424 552 486476 604
rect 489644 552 489696 604
rect 502984 552 503036 604
rect 446588 348 446640 400
rect 456708 348 456760 400
rect 453120 280 453172 332
rect 464160 280 464212 332
rect 237932 212 237984 264
rect 242256 212 242308 264
rect 353852 212 353904 264
rect 357348 212 357400 264
rect 390284 212 390336 264
rect 396356 212 396408 264
rect 401508 212 401560 264
rect 408592 212 408644 264
rect 412364 212 412416 264
rect 420368 212 420420 264
rect 423404 212 423456 264
rect 431868 212 431920 264
rect 434628 212 434680 264
rect 443644 212 443696 264
rect 445484 212 445536 264
rect 455880 212 455932 264
rect 456524 212 456576 264
rect 468852 484 468904 536
rect 480720 484 480772 536
rect 485412 484 485464 536
rect 498384 484 498436 536
rect 502800 484 502852 536
rect 517152 552 517204 604
rect 518440 552 518492 604
rect 519452 620 519504 672
rect 534816 620 534868 672
rect 529020 552 529072 604
rect 533712 552 533764 604
rect 535000 552 535052 604
rect 546684 688 546736 740
rect 536012 620 536064 672
rect 549076 552 549128 604
rect 506112 484 506164 536
rect 515772 484 515824 536
rect 551192 620 551244 672
rect 550272 552 550324 604
rect 550364 552 550416 604
rect 551376 688 551428 740
rect 569132 688 569184 740
rect 558092 620 558144 672
rect 576308 620 576360 672
rect 552664 552 552716 604
rect 479708 416 479760 468
rect 492496 416 492548 468
rect 496268 416 496320 468
rect 509884 416 509936 468
rect 512828 416 512880 468
rect 528008 416 528060 468
rect 529388 416 529440 468
rect 545672 416 545724 468
rect 568028 552 568080 604
rect 575112 552 575164 604
rect 556988 484 557040 536
rect 467656 348 467708 400
rect 479156 348 479208 400
rect 484216 348 484268 400
rect 497280 348 497332 400
rect 500776 348 500828 400
rect 514944 348 514996 400
rect 516140 348 516192 400
rect 531504 348 531556 400
rect 533896 348 533948 400
rect 549260 348 549312 400
rect 567016 416 567068 468
rect 555884 348 555936 400
rect 573732 348 573784 400
rect 473084 280 473136 332
rect 485044 280 485096 332
rect 485504 280 485556 332
rect 495716 280 495768 332
rect 499580 280 499632 332
rect 513380 280 513432 332
rect 522764 280 522816 332
rect 538220 280 538272 332
rect 539324 280 539376 332
rect 556344 280 556396 332
rect 556436 280 556488 332
rect 558736 280 558788 332
rect 560208 280 560260 332
rect 578792 280 578844 332
rect 471888 212 471940 264
rect 483848 212 483900 264
rect 488448 212 488500 264
rect 501604 212 501656 264
rect 505008 212 505060 264
rect 519728 212 519780 264
rect 521568 212 521620 264
rect 537392 212 537444 264
rect 538128 212 538180 264
rect 554780 212 554832 264
rect 563612 212 563664 264
rect 583576 212 583628 264
rect 223488 144 223540 196
rect 381452 144 381504 196
rect 386972 144 387024 196
rect 399944 144 399996 196
rect 407028 144 407080 196
rect 411168 144 411220 196
rect 418804 144 418856 196
rect 422208 144 422260 196
rect 431040 144 431092 196
rect 433064 144 433116 196
rect 442816 144 442868 196
rect 444288 144 444340 196
rect 454316 144 454368 196
rect 455328 144 455380 196
rect 466092 144 466144 196
rect 466460 144 466512 196
rect 478328 144 478380 196
rect 488632 144 488684 196
rect 490932 144 490984 196
rect 495164 144 495216 196
rect 509056 144 509108 196
rect 511724 144 511776 196
rect 526444 144 526496 196
rect 528284 144 528336 196
rect 544568 144 544620 196
rect 544844 144 544896 196
rect 562232 144 562284 196
rect 562508 144 562560 196
rect 582012 144 582064 196
rect 388 76 440 128
rect 20352 76 20404 128
rect 19616 8 19668 60
rect 38016 76 38068 128
rect 38568 76 38620 128
rect 55680 76 55732 128
rect 57060 76 57112 128
rect 73344 76 73396 128
rect 75184 76 75236 128
rect 89904 76 89956 128
rect 90180 76 90232 128
rect 104256 76 104308 128
rect 104348 76 104400 128
rect 117412 76 117464 128
rect 120908 76 120960 128
rect 132776 76 132828 128
rect 134340 76 134392 128
rect 145104 76 145156 128
rect 147312 8 147364 60
rect 157248 76 157300 128
rect 157984 76 158036 128
rect 167368 76 167420 128
rect 168656 76 168708 128
rect 177120 76 177172 128
rect 180432 76 180484 128
rect 188160 76 188212 128
rect 228548 76 228600 128
rect 232504 76 232556 128
rect 344928 76 344980 128
rect 348240 76 348292 128
rect 372528 76 372580 128
rect 377864 76 377916 128
rect 383384 76 383436 128
rect 389640 76 389692 128
rect 405648 76 405700 128
rect 412916 76 412968 128
rect 413468 76 413520 128
rect 421196 76 421248 128
rect 427728 76 427780 128
rect 436928 76 436980 128
rect 438768 76 438820 128
rect 448428 76 448480 128
rect 449624 76 449676 128
rect 460204 76 460256 128
rect 460848 76 460900 128
rect 472440 76 472492 128
rect 477408 76 477460 128
rect 490104 76 490156 128
rect 493968 76 494020 128
rect 507492 76 507544 128
rect 510528 76 510580 128
rect 525616 76 525668 128
rect 527088 76 527140 128
rect 543004 76 543056 128
rect 543648 76 543700 128
rect 560668 76 560720 128
rect 561404 76 561456 128
rect 581184 76 581236 128
rect 152004 8 152056 60
rect 161664 8 161716 60
rect 467288 8 467340 60
rect 470048 8 470100 60
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 20410 2802 20438 3060
rect 21514 2802 21542 3060
rect 22618 2802 22646 3060
rect 23722 2802 23750 3060
rect 24826 2802 24854 3060
rect 25930 2802 25958 3060
rect 27034 2802 27062 3060
rect 28138 2802 28166 3060
rect 29242 2802 29270 3060
rect 30346 2802 30374 3060
rect 31450 2802 31478 3060
rect 32554 2802 32582 3060
rect 33658 2802 33686 3060
rect 34762 2802 34790 3060
rect 35866 2802 35894 3060
rect 36970 2802 36998 3060
rect 38074 2802 38102 3060
rect 39178 2802 39206 3060
rect 40282 2802 40310 3060
rect 41386 2802 41414 3060
rect 42490 2802 42518 3060
rect 43594 2802 43622 3060
rect 44698 2802 44726 3060
rect 45802 2802 45830 3060
rect 46906 2802 46934 3060
rect 48010 2802 48038 3060
rect 20364 2774 20438 2802
rect 21468 2774 21542 2802
rect 22572 2774 22646 2802
rect 23676 2774 23750 2802
rect 24780 2774 24854 2802
rect 25884 2774 25958 2802
rect 26988 2774 27062 2802
rect 28092 2774 28166 2802
rect 29196 2774 29270 2802
rect 30300 2774 30374 2802
rect 31404 2774 31478 2802
rect 32508 2774 32582 2802
rect 33428 2774 33686 2802
rect 34532 2774 34790 2802
rect 35820 2774 35894 2802
rect 36924 2774 36998 2802
rect 38028 2774 38102 2802
rect 39132 2774 39206 2802
rect 40236 2774 40310 2802
rect 41340 2774 41414 2802
rect 42444 2774 42518 2802
rect 43548 2774 43622 2802
rect 44652 2774 44726 2802
rect 45756 2774 45830 2802
rect 46860 2774 46934 2802
rect 47964 2774 48038 2802
rect 49114 2802 49142 3060
rect 50218 2802 50246 3060
rect 51322 2802 51350 3060
rect 52426 2802 52454 3060
rect 53530 2802 53558 3060
rect 54634 2802 54662 3060
rect 55738 2802 55766 3060
rect 56842 2802 56870 3060
rect 57946 2802 57974 3060
rect 59050 2802 59078 3060
rect 59176 2916 59228 2922
rect 59176 2858 59228 2864
rect 49114 2774 49188 2802
rect 17040 1148 17092 1154
rect 17040 1090 17092 1096
rect 11152 876 11204 882
rect 11152 818 11204 824
rect 5264 672 5316 678
rect 5264 614 5316 620
rect 3882 504 3938 513
rect 388 128 440 134
rect 542 82 654 480
rect 1492 264 1544 270
rect 1646 218 1758 480
rect 1544 212 1758 218
rect 1492 206 1758 212
rect 1504 190 1758 206
rect 440 76 654 82
rect 388 70 654 76
rect 400 54 654 70
rect 542 -960 654 54
rect 1646 -960 1758 190
rect 2842 218 2954 480
rect 5276 480 5304 614
rect 6460 604 6512 610
rect 6460 546 6512 552
rect 6472 480 6500 546
rect 11164 480 11192 818
rect 12348 808 12400 814
rect 12348 750 12400 756
rect 12360 480 12388 750
rect 13544 740 13596 746
rect 13544 682 13596 688
rect 13556 480 13584 682
rect 14556 536 14608 542
rect 3882 439 3938 448
rect 3896 354 3924 439
rect 4038 354 4150 480
rect 3896 326 4150 354
rect 2842 202 3096 218
rect 2842 196 3108 202
rect 2842 190 3056 196
rect 2842 -960 2954 190
rect 3056 138 3108 144
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 354 7738 480
rect 7840 468 7892 474
rect 7840 410 7892 416
rect 7852 354 7880 410
rect 7626 326 7880 354
rect 8730 354 8842 480
rect 8944 400 8996 406
rect 8730 348 8944 354
rect 9926 354 10038 480
rect 8730 342 8996 348
rect 8730 326 8984 342
rect 9784 338 10038 354
rect 9772 332 10038 338
rect 7626 -960 7738 326
rect 8730 -960 8842 326
rect 9824 326 10038 332
rect 9772 274 9824 280
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14556 478 14608 484
rect 17052 480 17080 1090
rect 18236 1080 18288 1086
rect 18236 1022 18288 1028
rect 18248 480 18276 1022
rect 18880 1012 18932 1018
rect 18880 954 18932 960
rect 14568 354 14596 478
rect 14710 354 14822 480
rect 14568 326 14822 354
rect 14710 -960 14822 326
rect 15906 82 16018 480
rect 16210 96 16266 105
rect 15906 54 16210 82
rect 15906 -960 16018 54
rect 16210 31 16266 40
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 18892 202 18920 954
rect 18880 196 18932 202
rect 18880 138 18932 144
rect 19402 82 19514 480
rect 20364 134 20392 2774
rect 21180 944 21232 950
rect 21180 886 21232 892
rect 21192 610 21220 886
rect 21180 604 21232 610
rect 21180 546 21232 552
rect 20442 368 20498 377
rect 20598 354 20710 480
rect 21364 400 21416 406
rect 20498 326 20710 354
rect 21192 348 21364 354
rect 21192 342 21416 348
rect 21192 338 21404 342
rect 20442 303 20498 312
rect 20352 128 20404 134
rect 19402 66 19656 82
rect 20352 70 20404 76
rect 19402 60 19668 66
rect 19402 54 19616 60
rect 19402 -960 19514 54
rect 19616 2 19668 8
rect 20598 -960 20710 326
rect 21180 332 21404 338
rect 21232 326 21404 332
rect 21180 274 21232 280
rect 21468 202 21496 2774
rect 22572 1018 22600 2774
rect 23020 1284 23072 1290
rect 23020 1226 23072 1232
rect 22560 1012 22612 1018
rect 22560 954 22612 960
rect 23032 480 23060 1226
rect 23676 513 23704 2774
rect 24780 678 24808 2774
rect 25884 950 25912 2774
rect 25872 944 25924 950
rect 25872 886 25924 892
rect 24768 672 24820 678
rect 24768 614 24820 620
rect 24216 604 24268 610
rect 24216 546 24268 552
rect 25320 604 25372 610
rect 25320 546 25372 552
rect 23662 504 23718 513
rect 21794 218 21906 480
rect 22006 232 22062 241
rect 21456 196 21508 202
rect 21456 138 21508 144
rect 21794 190 22006 218
rect 21794 -960 21906 190
rect 22006 167 22062 176
rect 22990 -960 23102 480
rect 24228 480 24256 546
rect 25332 480 25360 546
rect 23662 439 23718 448
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26332 400 26384 406
rect 26486 354 26598 480
rect 26988 474 27016 2774
rect 26976 468 27028 474
rect 26976 410 27028 416
rect 26384 348 26598 354
rect 26332 342 26598 348
rect 26344 326 26598 342
rect 26486 -960 26598 326
rect 27682 218 27794 480
rect 28092 270 28120 2774
rect 28908 1352 28960 1358
rect 28908 1294 28960 1300
rect 28920 480 28948 1294
rect 28080 264 28132 270
rect 27682 202 27936 218
rect 28080 206 28132 212
rect 27682 196 27948 202
rect 27682 190 27896 196
rect 27682 -960 27794 190
rect 27896 138 27948 144
rect 28878 -960 28990 480
rect 29196 338 29224 2774
rect 30300 882 30328 2774
rect 30288 876 30340 882
rect 30288 818 30340 824
rect 30380 876 30432 882
rect 30380 818 30432 824
rect 30074 354 30186 480
rect 30392 354 30420 818
rect 31404 814 31432 2774
rect 31484 1216 31536 1222
rect 31484 1158 31536 1164
rect 31392 808 31444 814
rect 31392 750 31444 756
rect 31116 468 31168 474
rect 31116 410 31168 416
rect 29184 332 29236 338
rect 29184 274 29236 280
rect 30074 326 30420 354
rect 31128 354 31156 410
rect 31270 354 31382 480
rect 31496 406 31524 1158
rect 32508 746 32536 2774
rect 32496 740 32548 746
rect 32496 682 32548 688
rect 33428 542 33456 2774
rect 33612 598 33824 626
rect 33416 536 33468 542
rect 31128 326 31382 354
rect 31484 400 31536 406
rect 31484 342 31536 348
rect 32220 400 32272 406
rect 32374 354 32486 480
rect 33416 478 33468 484
rect 33612 480 33640 598
rect 32272 348 32486 354
rect 32220 342 32486 348
rect 32232 326 32486 342
rect 30074 -960 30186 326
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 33796 338 33824 598
rect 33784 332 33836 338
rect 33784 274 33836 280
rect 34426 96 34482 105
rect 34532 82 34560 2774
rect 35820 1018 35848 2774
rect 35992 1284 36044 1290
rect 35992 1226 36044 1232
rect 35808 1012 35860 1018
rect 35808 954 35860 960
rect 34796 808 34848 814
rect 34796 750 34848 756
rect 34808 480 34836 750
rect 36004 480 36032 1226
rect 36924 950 36952 2774
rect 36912 944 36964 950
rect 36912 886 36964 892
rect 37004 536 37056 542
rect 34482 54 34560 82
rect 34426 31 34482 40
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37004 478 37056 484
rect 37016 354 37044 478
rect 37158 354 37270 480
rect 37016 326 37270 354
rect 37158 -960 37270 326
rect 38028 134 38056 2774
rect 38016 128 38068 134
rect 38016 70 38068 76
rect 38354 82 38466 480
rect 39132 377 39160 2774
rect 39118 368 39174 377
rect 39118 303 39174 312
rect 38568 128 38620 134
rect 38354 76 38568 82
rect 38354 70 38620 76
rect 39394 96 39450 105
rect 38354 54 38608 70
rect 38354 -960 38466 54
rect 39550 82 39662 480
rect 40236 241 40264 2774
rect 41340 1086 41368 2774
rect 41328 1080 41380 1086
rect 41328 1022 41380 1028
rect 40684 1012 40736 1018
rect 40684 954 40736 960
rect 40696 480 40724 954
rect 41880 740 41932 746
rect 41880 682 41932 688
rect 41892 480 41920 682
rect 42444 678 42472 2774
rect 43548 678 43576 2774
rect 44652 1222 44680 2774
rect 44640 1216 44692 1222
rect 44640 1158 44692 1164
rect 42432 672 42484 678
rect 42432 614 42484 620
rect 43536 672 43588 678
rect 43536 614 43588 620
rect 43076 604 43128 610
rect 43076 546 43128 552
rect 43088 480 43116 546
rect 40222 232 40278 241
rect 40222 167 40278 176
rect 39450 54 39662 82
rect 39394 31 39450 40
rect 39550 -960 39662 54
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 218 44354 480
rect 44456 264 44508 270
rect 44242 212 44456 218
rect 44242 206 44508 212
rect 45282 232 45338 241
rect 44242 190 44496 206
rect 44242 -960 44354 190
rect 45438 218 45550 480
rect 45338 190 45550 218
rect 45756 202 45784 2774
rect 46860 1154 46888 2774
rect 46848 1148 46900 1154
rect 46848 1090 46900 1096
rect 46664 1080 46716 1086
rect 46664 1022 46716 1028
rect 46676 480 46704 1022
rect 47216 1012 47268 1018
rect 47216 954 47268 960
rect 47228 542 47256 954
rect 47964 882 47992 2774
rect 47952 876 48004 882
rect 47952 818 48004 824
rect 47860 740 47912 746
rect 47860 682 47912 688
rect 47216 536 47268 542
rect 45282 167 45338 176
rect 45438 -960 45550 190
rect 45744 196 45796 202
rect 45744 138 45796 144
rect 46634 -960 46746 480
rect 47216 478 47268 484
rect 47872 480 47900 682
rect 49160 542 49188 2774
rect 49988 2774 50246 2802
rect 51184 2774 51350 2802
rect 52380 2774 52454 2802
rect 53484 2774 53558 2802
rect 54588 2774 54662 2802
rect 55692 2774 55766 2802
rect 56796 2774 56870 2802
rect 57900 2774 57974 2802
rect 59004 2774 59078 2802
rect 49148 536 49200 542
rect 47830 -960 47942 480
rect 48780 468 48832 474
rect 48780 410 48832 416
rect 48792 354 48820 410
rect 48934 354 49046 480
rect 49148 478 49200 484
rect 49988 406 50016 2774
rect 50172 598 50384 626
rect 50172 480 50200 598
rect 48792 326 49046 354
rect 49976 400 50028 406
rect 49976 342 50028 348
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 50356 202 50384 598
rect 51184 338 51212 2774
rect 51356 1216 51408 1222
rect 51356 1158 51408 1164
rect 51368 480 51396 1158
rect 52380 814 52408 2774
rect 53484 1290 53512 2774
rect 53472 1284 53524 1290
rect 53472 1226 53524 1232
rect 54588 1018 54616 2774
rect 54576 1012 54628 1018
rect 54576 954 54628 960
rect 52368 808 52420 814
rect 52368 750 52420 756
rect 53748 808 53800 814
rect 53748 750 53800 756
rect 52552 740 52604 746
rect 52552 682 52604 688
rect 52564 480 52592 682
rect 53760 480 53788 750
rect 51172 332 51224 338
rect 51172 274 51224 280
rect 50344 196 50396 202
rect 50344 138 50396 144
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 354 55026 480
rect 55128 400 55180 406
rect 54914 348 55128 354
rect 54914 342 55180 348
rect 54914 326 55168 342
rect 54914 -960 55026 326
rect 55692 134 55720 2774
rect 56018 354 56130 480
rect 56018 338 56272 354
rect 56018 332 56284 338
rect 56018 326 56232 332
rect 55680 128 55732 134
rect 55680 70 55732 76
rect 56018 -960 56130 326
rect 56232 274 56284 280
rect 56796 105 56824 2774
rect 57900 950 57928 2774
rect 58440 1148 58492 1154
rect 58440 1090 58492 1096
rect 57888 944 57940 950
rect 57888 886 57940 892
rect 58452 480 58480 1090
rect 59004 678 59032 2774
rect 59188 882 59216 2858
rect 60154 2802 60182 3060
rect 61258 2802 61286 3060
rect 60108 2774 60182 2802
rect 61212 2774 61286 2802
rect 62362 2802 62390 3060
rect 63466 2938 63494 3060
rect 63420 2910 63494 2938
rect 64570 2922 64598 3060
rect 64558 2916 64610 2922
rect 62362 2774 62436 2802
rect 59636 944 59688 950
rect 59636 886 59688 892
rect 59176 876 59228 882
rect 59176 818 59228 824
rect 58992 672 59044 678
rect 58992 614 59044 620
rect 59648 480 59676 886
rect 60108 610 60136 2774
rect 60832 876 60884 882
rect 60832 818 60884 824
rect 60096 604 60148 610
rect 60096 546 60148 552
rect 60844 480 60872 818
rect 57060 128 57112 134
rect 56782 96 56838 105
rect 57214 82 57326 480
rect 57112 76 57326 82
rect 57060 70 57326 76
rect 57072 54 57326 70
rect 56782 31 56838 40
rect 57214 -960 57326 54
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61212 270 61240 2774
rect 62028 604 62080 610
rect 62028 546 62080 552
rect 62040 480 62068 546
rect 61200 264 61252 270
rect 61200 206 61252 212
rect 61998 -960 62110 480
rect 62408 241 62436 2774
rect 63420 1018 63448 2910
rect 64558 2858 64610 2864
rect 63500 2848 63552 2854
rect 63500 2790 63552 2796
rect 65674 2802 65702 3060
rect 66778 2802 66806 3060
rect 67640 2916 67692 2922
rect 67640 2858 67692 2864
rect 63512 1086 63540 2790
rect 65674 2774 65748 2802
rect 65524 1216 65576 1222
rect 65524 1158 65576 1164
rect 63500 1080 63552 1086
rect 63500 1022 63552 1028
rect 63408 1012 63460 1018
rect 63408 954 63460 960
rect 64328 672 64380 678
rect 64328 614 64380 620
rect 64340 480 64368 614
rect 65536 480 65564 1158
rect 62394 232 62450 241
rect 62394 167 62450 176
rect 63194 218 63306 480
rect 63408 264 63460 270
rect 63194 212 63408 218
rect 63194 206 63460 212
rect 63194 190 63448 206
rect 63194 -960 63306 190
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 65720 474 65748 2774
rect 66548 2774 66806 2802
rect 65708 468 65760 474
rect 65708 410 65760 416
rect 66548 202 66576 2774
rect 67652 814 67680 2858
rect 67882 2854 67910 3060
rect 67870 2848 67922 2854
rect 68986 2802 69014 3060
rect 70090 2922 70118 3060
rect 70078 2916 70130 2922
rect 70078 2858 70130 2864
rect 71194 2802 71222 3060
rect 71780 2916 71832 2922
rect 71780 2858 71832 2864
rect 67870 2790 67922 2796
rect 68940 2774 69014 2802
rect 71148 2774 71222 2802
rect 67640 808 67692 814
rect 67640 750 67692 756
rect 68940 746 68968 2774
rect 69112 1080 69164 1086
rect 69112 1022 69164 1028
rect 68928 740 68980 746
rect 68928 682 68980 688
rect 67928 598 68140 626
rect 66732 564 66944 592
rect 66732 480 66760 564
rect 66536 196 66588 202
rect 66536 138 66588 144
rect 66690 -960 66802 480
rect 66916 474 66944 564
rect 67928 480 67956 598
rect 66904 468 66956 474
rect 66904 410 66956 416
rect 67886 -960 67998 480
rect 68112 354 68140 598
rect 69124 480 69152 1022
rect 70308 740 70360 746
rect 70308 682 70360 688
rect 70320 480 70348 682
rect 68112 326 68232 354
rect 68204 202 68232 326
rect 68192 196 68244 202
rect 68192 138 68244 144
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71148 406 71176 2774
rect 71792 1154 71820 2858
rect 72298 2802 72326 3060
rect 72252 2774 72326 2802
rect 73160 2848 73212 2854
rect 73402 2802 73430 3060
rect 74506 2922 74534 3060
rect 74494 2916 74546 2922
rect 74494 2858 74546 2864
rect 75460 2916 75512 2922
rect 75460 2858 75512 2864
rect 73160 2790 73212 2796
rect 71780 1148 71832 1154
rect 71780 1090 71832 1096
rect 71504 1012 71556 1018
rect 71504 954 71556 960
rect 71516 480 71544 954
rect 71136 400 71188 406
rect 71136 342 71188 348
rect 71474 -960 71586 480
rect 72252 338 72280 2774
rect 73172 950 73200 2790
rect 73356 2774 73430 2802
rect 73160 944 73212 950
rect 73160 886 73212 892
rect 72608 808 72660 814
rect 72608 750 72660 756
rect 72620 480 72648 750
rect 72240 332 72292 338
rect 72240 274 72292 280
rect 72578 -960 72690 480
rect 73356 134 73384 2774
rect 75472 678 75500 2858
rect 75610 2854 75638 3060
rect 76714 2922 76742 3060
rect 76702 2916 76754 2922
rect 76702 2858 76754 2864
rect 75598 2848 75650 2854
rect 75598 2790 75650 2796
rect 76840 2848 76892 2854
rect 77818 2802 77846 3060
rect 78922 2802 78950 3060
rect 80026 2938 80054 3060
rect 76840 2790 76892 2796
rect 76852 1154 76880 2790
rect 77772 2774 77846 2802
rect 78876 2774 78950 2802
rect 79980 2910 80054 2938
rect 80152 2916 80204 2922
rect 76840 1148 76892 1154
rect 76840 1090 76892 1096
rect 77392 1148 77444 1154
rect 77392 1090 77444 1096
rect 76932 876 76984 882
rect 76932 818 76984 824
rect 75460 672 75512 678
rect 75460 614 75512 620
rect 76196 672 76248 678
rect 76196 614 76248 620
rect 76208 480 76236 614
rect 73774 354 73886 480
rect 73632 338 73886 354
rect 73620 332 73886 338
rect 73672 326 73886 332
rect 73620 274 73672 280
rect 73344 128 73396 134
rect 73344 70 73396 76
rect 73774 -960 73886 326
rect 74970 82 75082 480
rect 75184 128 75236 134
rect 74970 76 75184 82
rect 74970 70 75236 76
rect 74970 54 75224 70
rect 74970 -960 75082 54
rect 76166 -960 76278 480
rect 76944 474 76972 818
rect 77404 480 77432 1090
rect 77772 542 77800 2774
rect 77760 536 77812 542
rect 76932 468 76984 474
rect 76932 410 76984 416
rect 77362 -960 77474 480
rect 77760 478 77812 484
rect 78404 400 78456 406
rect 78558 354 78670 480
rect 78456 348 78670 354
rect 78404 342 78670 348
rect 78416 326 78670 342
rect 78558 -960 78670 326
rect 78876 270 78904 2774
rect 79692 604 79744 610
rect 79692 546 79744 552
rect 79704 480 79732 546
rect 78864 264 78916 270
rect 78864 206 78916 212
rect 79662 -960 79774 480
rect 79980 474 80008 2910
rect 80152 2858 80204 2864
rect 80164 1086 80192 2858
rect 81130 2854 81158 3060
rect 81118 2848 81170 2854
rect 82234 2802 82262 3060
rect 83338 2802 83366 3060
rect 84442 2922 84470 3060
rect 84430 2916 84482 2922
rect 84430 2858 84482 2864
rect 85396 2916 85448 2922
rect 85396 2858 85448 2864
rect 81118 2790 81170 2796
rect 82188 2774 82262 2802
rect 83108 2774 83366 2802
rect 80152 1080 80204 1086
rect 80152 1022 80204 1028
rect 82188 882 82216 2774
rect 82176 876 82228 882
rect 82176 818 82228 824
rect 82084 604 82136 610
rect 82084 546 82136 552
rect 82096 480 82124 546
rect 79968 468 80020 474
rect 79968 410 80020 416
rect 80858 218 80970 480
rect 81072 264 81124 270
rect 80858 212 81072 218
rect 80858 206 81124 212
rect 80858 190 81112 206
rect 80858 -960 80970 190
rect 82054 -960 82166 480
rect 83108 202 83136 2774
rect 85408 1018 85436 2858
rect 85546 2802 85574 3060
rect 86650 2922 86678 3060
rect 87754 2922 87782 3060
rect 86638 2916 86690 2922
rect 86638 2858 86690 2864
rect 86776 2916 86828 2922
rect 86776 2858 86828 2864
rect 87742 2916 87794 2922
rect 87742 2858 87794 2864
rect 88156 2916 88208 2922
rect 88156 2858 88208 2864
rect 85500 2774 85574 2802
rect 85396 1012 85448 1018
rect 85396 954 85448 960
rect 83280 944 83332 950
rect 83280 886 83332 892
rect 83292 480 83320 886
rect 85500 746 85528 2774
rect 86788 814 86816 2858
rect 88168 1154 88196 2858
rect 88858 2802 88886 3060
rect 89962 2802 89990 3060
rect 91066 2802 91094 3060
rect 92170 2922 92198 3060
rect 92158 2916 92210 2922
rect 92158 2858 92210 2864
rect 92480 2916 92532 2922
rect 92480 2858 92532 2864
rect 88812 2774 88886 2802
rect 89916 2774 89990 2802
rect 91020 2774 91094 2802
rect 88156 1148 88208 1154
rect 88156 1090 88208 1096
rect 86868 944 86920 950
rect 86868 886 86920 892
rect 86776 808 86828 814
rect 86776 750 86828 756
rect 85488 740 85540 746
rect 85488 682 85540 688
rect 84488 598 84700 626
rect 84488 480 84516 598
rect 83096 196 83148 202
rect 83096 138 83148 144
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 84672 474 84700 598
rect 86880 480 86908 886
rect 87972 740 88024 746
rect 87972 682 88024 688
rect 87984 480 88012 682
rect 84660 468 84712 474
rect 84660 410 84712 416
rect 85642 218 85754 480
rect 85642 202 85896 218
rect 85642 196 85908 202
rect 85642 190 85856 196
rect 85642 -960 85754 190
rect 85856 138 85908 144
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 88812 338 88840 2774
rect 89168 808 89220 814
rect 89168 750 89220 756
rect 89180 480 89208 750
rect 88800 332 88852 338
rect 88800 274 88852 280
rect 89138 -960 89250 480
rect 89916 134 89944 2774
rect 91020 678 91048 2774
rect 91560 1012 91612 1018
rect 91560 954 91612 960
rect 91008 672 91060 678
rect 91008 614 91060 620
rect 91572 480 91600 954
rect 92492 542 92520 2858
rect 93274 2802 93302 3060
rect 94378 2922 94406 3060
rect 95482 2922 95510 3060
rect 94366 2916 94418 2922
rect 94366 2858 94418 2864
rect 94596 2916 94648 2922
rect 94596 2858 94648 2864
rect 95470 2916 95522 2922
rect 95470 2858 95522 2864
rect 95700 2916 95752 2922
rect 95700 2858 95752 2864
rect 93228 2774 93302 2802
rect 92480 536 92532 542
rect 89904 128 89956 134
rect 89904 70 89956 76
rect 90180 128 90232 134
rect 90334 82 90446 480
rect 90232 76 90446 82
rect 90180 70 90446 76
rect 90192 54 90446 70
rect 90334 -960 90446 54
rect 91530 -960 91642 480
rect 92480 478 92532 484
rect 92572 400 92624 406
rect 92726 354 92838 480
rect 92624 348 92838 354
rect 92572 342 92838 348
rect 92584 326 92838 342
rect 93228 338 93256 2774
rect 93922 354 94034 480
rect 93922 338 94176 354
rect 92726 -960 92838 326
rect 93216 332 93268 338
rect 93216 274 93268 280
rect 93922 332 94188 338
rect 93922 326 94136 332
rect 93922 -960 94034 326
rect 94136 274 94188 280
rect 94608 270 94636 2858
rect 95712 882 95740 2858
rect 96586 2802 96614 3060
rect 97690 2922 97718 3060
rect 97678 2916 97730 2922
rect 97678 2858 97730 2864
rect 98000 2916 98052 2922
rect 98000 2858 98052 2864
rect 96540 2774 96614 2802
rect 95700 876 95752 882
rect 95700 818 95752 824
rect 96252 740 96304 746
rect 96252 682 96304 688
rect 95148 672 95200 678
rect 95148 614 95200 620
rect 95160 480 95188 614
rect 96264 480 96292 682
rect 96540 610 96568 2774
rect 97448 1080 97500 1086
rect 97448 1022 97500 1028
rect 96528 604 96580 610
rect 96528 546 96580 552
rect 97460 480 97488 1022
rect 98012 950 98040 2858
rect 98794 2802 98822 3060
rect 99898 2802 99926 3060
rect 101002 2922 101030 3060
rect 102106 2938 102134 3060
rect 100990 2916 101042 2922
rect 100990 2858 101042 2864
rect 102060 2910 102134 2938
rect 102232 2916 102284 2922
rect 98794 2774 98868 2802
rect 98000 944 98052 950
rect 98000 886 98052 892
rect 94596 264 94648 270
rect 94596 206 94648 212
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98460 264 98512 270
rect 98614 218 98726 480
rect 98840 474 98868 2774
rect 99668 2774 99926 2802
rect 100760 2848 100812 2854
rect 100760 2790 100812 2796
rect 98828 468 98880 474
rect 98828 410 98880 416
rect 98512 212 98726 218
rect 98460 206 98726 212
rect 98472 190 98726 206
rect 99668 202 99696 2774
rect 100772 950 100800 2790
rect 100760 944 100812 950
rect 100760 886 100812 892
rect 99840 876 99892 882
rect 99840 818 99892 824
rect 99852 480 99880 818
rect 102060 814 102088 2910
rect 102232 2858 102284 2864
rect 102244 1018 102272 2858
rect 103210 2854 103238 3060
rect 103198 2848 103250 2854
rect 104314 2802 104342 3060
rect 105418 2922 105446 3060
rect 106522 2922 106550 3060
rect 105406 2916 105458 2922
rect 105406 2858 105458 2864
rect 105544 2916 105596 2922
rect 105544 2858 105596 2864
rect 106510 2916 106562 2922
rect 106510 2858 106562 2864
rect 103198 2790 103250 2796
rect 104268 2774 104342 2802
rect 102232 1012 102284 1018
rect 102232 954 102284 960
rect 102048 808 102100 814
rect 102048 750 102100 756
rect 103336 740 103388 746
rect 103336 682 103388 688
rect 101312 672 101364 678
rect 101312 614 101364 620
rect 101036 604 101088 610
rect 101036 546 101088 552
rect 101048 480 101076 546
rect 98614 -960 98726 190
rect 99656 196 99708 202
rect 99656 138 99708 144
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 101324 338 101352 614
rect 103348 480 103376 682
rect 101312 332 101364 338
rect 101312 274 101364 280
rect 102202 218 102314 480
rect 102202 202 102456 218
rect 102202 196 102468 202
rect 102202 190 102416 196
rect 102202 -960 102314 190
rect 102416 138 102468 144
rect 103306 -960 103418 480
rect 104268 134 104296 2774
rect 104256 128 104308 134
rect 104256 70 104308 76
rect 104348 128 104400 134
rect 104502 82 104614 480
rect 105556 406 105584 2858
rect 107626 2802 107654 3060
rect 107752 2916 107804 2922
rect 107752 2858 107804 2864
rect 107580 2774 107654 2802
rect 105728 944 105780 950
rect 105728 886 105780 892
rect 105740 480 105768 886
rect 106004 808 106056 814
rect 106004 750 106056 756
rect 106016 610 106044 750
rect 107580 678 107608 2774
rect 107764 814 107792 2858
rect 108730 2802 108758 3060
rect 109834 2922 109862 3060
rect 109822 2916 109874 2922
rect 109822 2858 109874 2864
rect 110420 2916 110472 2922
rect 110420 2858 110472 2864
rect 108684 2774 108758 2802
rect 107752 808 107804 814
rect 107752 750 107804 756
rect 107568 672 107620 678
rect 107568 614 107620 620
rect 106004 604 106056 610
rect 106004 546 106056 552
rect 108120 604 108172 610
rect 108120 546 108172 552
rect 106740 536 106792 542
rect 105544 400 105596 406
rect 105544 342 105596 348
rect 104400 76 104614 82
rect 104348 70 104614 76
rect 104360 54 104614 70
rect 104502 -960 104614 54
rect 105698 -960 105810 480
rect 106740 478 106792 484
rect 108132 480 108160 546
rect 106752 354 106780 478
rect 106894 354 107006 480
rect 106752 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 108684 406 108712 2774
rect 110432 882 110460 2858
rect 110938 2802 110966 3060
rect 112042 2802 112070 3060
rect 113146 2922 113174 3060
rect 113134 2916 113186 2922
rect 113134 2858 113186 2864
rect 114250 2802 114278 3060
rect 114744 2916 114796 2922
rect 114744 2858 114796 2864
rect 110892 2774 110966 2802
rect 111996 2774 112070 2802
rect 114204 2774 114278 2802
rect 110892 1086 110920 2774
rect 110880 1080 110932 1086
rect 110880 1022 110932 1028
rect 111616 1080 111668 1086
rect 111616 1022 111668 1028
rect 110420 876 110472 882
rect 110420 818 110472 824
rect 111628 480 111656 1022
rect 108672 400 108724 406
rect 108672 342 108724 348
rect 109132 400 109184 406
rect 109286 354 109398 480
rect 109184 348 109398 354
rect 109132 342 109398 348
rect 109144 326 109398 342
rect 109286 -960 109398 326
rect 110482 354 110594 480
rect 110482 338 110736 354
rect 110482 332 110748 338
rect 110482 326 110696 332
rect 110482 -960 110594 326
rect 110696 274 110748 280
rect 111586 -960 111698 480
rect 111996 270 112024 2774
rect 112812 808 112864 814
rect 112812 750 112864 756
rect 112824 480 112852 750
rect 114204 542 114232 2774
rect 114756 1154 114784 2858
rect 115354 2802 115382 3060
rect 116458 2922 116486 3060
rect 116446 2916 116498 2922
rect 116446 2858 116498 2864
rect 117320 2916 117372 2922
rect 117320 2858 117372 2864
rect 115354 2774 115428 2802
rect 114744 1148 114796 1154
rect 114744 1090 114796 1096
rect 115204 876 115256 882
rect 115204 818 115256 824
rect 114192 536 114244 542
rect 111984 264 112036 270
rect 111984 206 112036 212
rect 112782 -960 112894 480
rect 113978 218 114090 480
rect 114192 478 114244 484
rect 115216 480 115244 818
rect 114192 264 114244 270
rect 113978 212 114192 218
rect 113978 206 114244 212
rect 113978 190 114232 206
rect 113978 -960 114090 190
rect 115174 -960 115286 480
rect 115400 202 115428 2774
rect 117332 950 117360 2858
rect 117562 2802 117590 3060
rect 118666 2802 118694 3060
rect 119770 2922 119798 3060
rect 119758 2916 119810 2922
rect 119758 2858 119810 2864
rect 120080 2916 120132 2922
rect 120080 2858 120132 2864
rect 117424 2774 117590 2802
rect 118620 2774 118694 2802
rect 117320 944 117372 950
rect 117320 886 117372 892
rect 116412 598 116624 626
rect 116412 480 116440 598
rect 115388 196 115440 202
rect 115388 138 115440 144
rect 116370 -960 116482 480
rect 116596 202 116624 598
rect 116584 196 116636 202
rect 116584 138 116636 144
rect 117424 134 117452 2774
rect 118620 1222 118648 2774
rect 118608 1216 118660 1222
rect 118608 1158 118660 1164
rect 120092 950 120120 2858
rect 120874 2802 120902 3060
rect 121978 2802 122006 3060
rect 123082 2802 123110 3060
rect 124186 2922 124214 3060
rect 124174 2916 124226 2922
rect 124174 2858 124226 2864
rect 125140 2916 125192 2922
rect 125140 2858 125192 2864
rect 120828 2774 120902 2802
rect 121932 2774 122006 2802
rect 123036 2774 123110 2802
rect 120080 944 120132 950
rect 120080 886 120132 892
rect 117596 740 117648 746
rect 117596 682 117648 688
rect 117608 480 117636 682
rect 118792 672 118844 678
rect 118792 614 118844 620
rect 118804 480 118832 614
rect 120828 542 120856 2774
rect 120816 536 120868 542
rect 117412 128 117464 134
rect 117412 70 117464 76
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 354 119978 480
rect 120816 478 120868 484
rect 120080 468 120132 474
rect 120080 410 120132 416
rect 120092 354 120120 410
rect 119866 326 120120 354
rect 119866 -960 119978 326
rect 120908 128 120960 134
rect 121062 82 121174 480
rect 121932 406 121960 2774
rect 121920 400 121972 406
rect 121920 342 121972 348
rect 122258 354 122370 480
rect 122472 400 122524 406
rect 122258 348 122472 354
rect 122258 342 122524 348
rect 120960 76 121174 82
rect 120908 70 121174 76
rect 120920 54 121174 70
rect 121062 -960 121174 54
rect 122258 326 122512 342
rect 123036 338 123064 2774
rect 125152 882 125180 2858
rect 125290 2802 125318 3060
rect 126394 2802 126422 3060
rect 127498 2922 127526 3060
rect 127486 2916 127538 2922
rect 127486 2858 127538 2864
rect 127624 2916 127676 2922
rect 127624 2858 127676 2864
rect 125244 2774 125318 2802
rect 126348 2774 126422 2802
rect 125140 876 125192 882
rect 125140 818 125192 824
rect 123484 808 123536 814
rect 123484 750 123536 756
rect 123496 480 123524 750
rect 125244 610 125272 2774
rect 125232 604 125284 610
rect 125232 546 125284 552
rect 124864 536 124916 542
rect 123024 332 123076 338
rect 122258 -960 122370 326
rect 123024 274 123076 280
rect 123454 -960 123566 480
rect 124650 354 124762 480
rect 124864 478 124916 484
rect 124876 354 124904 478
rect 125846 354 125958 480
rect 124650 326 124904 354
rect 125704 338 125958 354
rect 125692 332 125958 338
rect 124650 -960 124762 326
rect 125744 326 125958 332
rect 125692 274 125744 280
rect 125846 -960 125958 326
rect 126348 270 126376 2774
rect 127532 944 127584 950
rect 127532 886 127584 892
rect 126336 264 126388 270
rect 126336 206 126388 212
rect 126796 264 126848 270
rect 126950 218 127062 480
rect 127544 406 127572 886
rect 127636 746 127664 2858
rect 128602 2802 128630 3060
rect 129706 2922 129734 3060
rect 129694 2916 129746 2922
rect 129694 2858 129746 2864
rect 130810 2802 130838 3060
rect 128556 2774 128630 2802
rect 130764 2774 130838 2802
rect 131914 2802 131942 3060
rect 133018 2802 133046 3060
rect 134122 2922 134150 3060
rect 133236 2916 133288 2922
rect 133236 2858 133288 2864
rect 134110 2916 134162 2922
rect 134110 2858 134162 2864
rect 131914 2774 131988 2802
rect 128176 876 128228 882
rect 128176 818 128228 824
rect 127624 740 127676 746
rect 127624 682 127676 688
rect 128188 480 128216 818
rect 127532 400 127584 406
rect 127532 342 127584 348
rect 126848 212 127062 218
rect 126796 206 127062 212
rect 126808 190 127062 206
rect 126950 -960 127062 190
rect 128146 -960 128258 480
rect 128556 202 128584 2774
rect 129372 808 129424 814
rect 129372 750 129424 756
rect 129384 480 129412 750
rect 130764 678 130792 2774
rect 130752 672 130804 678
rect 130752 614 130804 620
rect 130568 604 130620 610
rect 130568 546 130620 552
rect 130580 480 130608 546
rect 128544 196 128596 202
rect 128544 138 128596 144
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131580 468 131632 474
rect 131580 410 131632 416
rect 131592 354 131620 410
rect 131734 354 131846 480
rect 131960 406 131988 2774
rect 132788 2774 133046 2802
rect 131592 326 131846 354
rect 131948 400 132000 406
rect 131948 342 132000 348
rect 131734 -960 131846 326
rect 132788 134 132816 2774
rect 133248 950 133276 2858
rect 135226 2802 135254 3060
rect 136330 2802 136358 3060
rect 136640 2916 136692 2922
rect 136640 2858 136692 2864
rect 135180 2774 135254 2802
rect 136284 2774 136358 2802
rect 133236 944 133288 950
rect 133236 886 133288 892
rect 135180 746 135208 2774
rect 135260 944 135312 950
rect 135260 886 135312 892
rect 135168 740 135220 746
rect 135168 682 135220 688
rect 132972 598 133184 626
rect 132972 480 133000 598
rect 132776 128 132828 134
rect 132776 70 132828 76
rect 132930 -960 133042 480
rect 133156 202 133184 598
rect 134168 598 134380 626
rect 134168 480 134196 598
rect 133144 196 133196 202
rect 133144 138 133196 144
rect 134126 -960 134238 480
rect 134352 134 134380 598
rect 135272 480 135300 886
rect 136284 542 136312 2774
rect 136652 882 136680 2858
rect 137434 2802 137462 3060
rect 138538 2802 138566 3060
rect 139642 2922 139670 3060
rect 139630 2916 139682 2922
rect 139630 2858 139682 2864
rect 140746 2802 140774 3060
rect 141850 2802 141878 3060
rect 142954 2802 142982 3060
rect 144058 2802 144086 3060
rect 144184 2916 144236 2922
rect 144184 2858 144236 2864
rect 137388 2774 137462 2802
rect 138492 2774 138566 2802
rect 140700 2774 140774 2802
rect 141804 2774 141878 2802
rect 142908 2774 142982 2802
rect 144012 2774 144086 2802
rect 136640 876 136692 882
rect 136640 818 136692 824
rect 136456 672 136508 678
rect 136456 614 136508 620
rect 136272 536 136324 542
rect 134340 128 134392 134
rect 134340 70 134392 76
rect 135230 -960 135342 480
rect 136272 478 136324 484
rect 136468 480 136496 614
rect 136426 -960 136538 480
rect 137388 338 137416 2774
rect 137468 400 137520 406
rect 137622 354 137734 480
rect 137520 348 137734 354
rect 137468 342 137734 348
rect 137376 332 137428 338
rect 137480 326 137734 342
rect 137376 274 137428 280
rect 137622 -960 137734 326
rect 138492 270 138520 2774
rect 140044 876 140096 882
rect 140044 818 140096 824
rect 140056 480 140084 818
rect 140700 814 140728 2774
rect 140688 808 140740 814
rect 140688 750 140740 756
rect 141240 808 141292 814
rect 141240 750 141292 756
rect 141252 480 141280 750
rect 141804 610 141832 2774
rect 141792 604 141844 610
rect 141792 546 141844 552
rect 142436 604 142488 610
rect 142436 546 142488 552
rect 142448 480 142476 546
rect 138818 354 138930 480
rect 138818 338 139072 354
rect 138818 332 139084 338
rect 138818 326 139032 332
rect 138480 264 138532 270
rect 138480 206 138532 212
rect 138818 -960 138930 326
rect 139032 274 139084 280
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 142908 474 142936 2774
rect 143448 1012 143500 1018
rect 143448 954 143500 960
rect 143460 814 143488 954
rect 143448 808 143500 814
rect 143448 750 143500 756
rect 143540 808 143592 814
rect 143540 750 143592 756
rect 143552 480 143580 750
rect 142896 468 142948 474
rect 142896 410 142948 416
rect 143510 -960 143622 480
rect 144012 202 144040 2774
rect 144196 950 144224 2858
rect 145162 2802 145190 3060
rect 146266 2922 146294 3060
rect 146254 2916 146306 2922
rect 146254 2858 146306 2864
rect 147370 2802 147398 3060
rect 145116 2774 145190 2802
rect 147324 2774 147398 2802
rect 148474 2802 148502 3060
rect 149060 2916 149112 2922
rect 149060 2858 149112 2864
rect 148474 2774 148548 2802
rect 144184 944 144236 950
rect 144184 886 144236 892
rect 144736 740 144788 746
rect 144736 682 144788 688
rect 144748 480 144776 682
rect 144000 196 144052 202
rect 144000 138 144052 144
rect 144706 -960 144818 480
rect 145116 134 145144 2774
rect 147324 678 147352 2774
rect 148324 944 148376 950
rect 148324 886 148376 892
rect 147312 672 147364 678
rect 147312 614 147364 620
rect 148336 480 148364 886
rect 145748 468 145800 474
rect 145748 410 145800 416
rect 145760 354 145788 410
rect 145902 354 146014 480
rect 145760 326 146014 354
rect 145104 128 145156 134
rect 145104 70 145156 76
rect 145902 -960 146014 326
rect 147098 82 147210 480
rect 147098 66 147352 82
rect 147098 60 147364 66
rect 147098 54 147312 60
rect 147098 -960 147210 54
rect 147312 2 147364 8
rect 148294 -960 148406 480
rect 148520 406 148548 2774
rect 149072 1018 149100 2858
rect 149578 2802 149606 3060
rect 149348 2774 149606 2802
rect 150440 2848 150492 2854
rect 150682 2802 150710 3060
rect 151786 2922 151814 3060
rect 151774 2916 151826 2922
rect 151774 2858 151826 2864
rect 152890 2854 152918 3060
rect 153384 2916 153436 2922
rect 153384 2858 153436 2864
rect 150440 2790 150492 2796
rect 149060 1012 149112 1018
rect 149060 954 149112 960
rect 148508 400 148560 406
rect 148508 342 148560 348
rect 149348 338 149376 2774
rect 149520 672 149572 678
rect 149520 614 149572 620
rect 149532 480 149560 614
rect 150452 610 150480 2790
rect 150636 2774 150710 2802
rect 152878 2848 152930 2854
rect 152878 2790 152930 2796
rect 150636 882 150664 2774
rect 150624 876 150676 882
rect 150624 818 150676 824
rect 153396 746 153424 2858
rect 153994 2802 154022 3060
rect 155098 2922 155126 3060
rect 155086 2916 155138 2922
rect 155086 2858 155138 2864
rect 155960 2916 156012 2922
rect 155960 2858 156012 2864
rect 153948 2774 154022 2802
rect 153948 814 153976 2774
rect 155972 950 156000 2858
rect 156202 2802 156230 3060
rect 157306 2802 157334 3060
rect 158410 2922 158438 3060
rect 158398 2916 158450 2922
rect 158398 2858 158450 2864
rect 158720 2916 158772 2922
rect 158720 2858 158772 2864
rect 156156 2774 156230 2802
rect 157260 2774 157334 2802
rect 155960 944 156012 950
rect 155960 886 156012 892
rect 153936 808 153988 814
rect 153936 750 153988 756
rect 153384 740 153436 746
rect 153384 682 153436 688
rect 150440 604 150492 610
rect 150440 546 150492 552
rect 150624 604 150676 610
rect 150624 546 150676 552
rect 151832 598 152044 626
rect 150636 480 150664 546
rect 151832 480 151860 598
rect 149336 332 149388 338
rect 149336 274 149388 280
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152016 66 152044 598
rect 154212 604 154264 610
rect 154212 546 154264 552
rect 154224 480 154252 546
rect 152986 354 153098 480
rect 152986 338 153240 354
rect 152986 332 153252 338
rect 152986 326 153200 332
rect 152004 60 152056 66
rect 152004 2 152056 8
rect 152986 -960 153098 326
rect 153200 274 153252 280
rect 154182 -960 154294 480
rect 155378 354 155490 480
rect 155592 400 155644 406
rect 155378 348 155592 354
rect 155378 342 155644 348
rect 155378 326 155632 342
rect 155378 -960 155490 326
rect 156156 202 156184 2774
rect 156420 468 156472 474
rect 156420 410 156472 416
rect 156432 354 156460 410
rect 156574 354 156686 480
rect 156432 326 156686 354
rect 156144 196 156196 202
rect 156144 138 156196 144
rect 156574 -960 156686 326
rect 157260 134 157288 2774
rect 157248 128 157300 134
rect 157248 70 157300 76
rect 157770 82 157882 480
rect 158732 338 158760 2858
rect 159514 2802 159542 3060
rect 160618 2802 160646 3060
rect 161722 2802 161750 3060
rect 162826 2922 162854 3060
rect 162814 2916 162866 2922
rect 162814 2858 162866 2864
rect 163930 2802 163958 3060
rect 159468 2774 159542 2802
rect 160572 2774 160646 2802
rect 161676 2774 161750 2802
rect 163884 2774 163958 2802
rect 165034 2802 165062 3060
rect 166138 2802 166166 3060
rect 167000 2916 167052 2922
rect 167000 2858 167052 2864
rect 165034 2774 165108 2802
rect 159468 678 159496 2774
rect 159456 672 159508 678
rect 159456 614 159508 620
rect 160100 672 160152 678
rect 160100 614 160152 620
rect 160112 480 160140 614
rect 158874 354 158986 480
rect 158874 338 159128 354
rect 158720 332 158772 338
rect 158720 274 158772 280
rect 158874 332 159140 338
rect 158874 326 159088 332
rect 157984 128 158036 134
rect 157770 76 157984 82
rect 157770 70 158036 76
rect 157770 54 158024 70
rect 157770 -960 157882 54
rect 158874 -960 158986 326
rect 159088 274 159140 280
rect 160070 -960 160182 480
rect 160572 270 160600 2774
rect 161480 876 161532 882
rect 161480 818 161532 824
rect 161266 354 161378 480
rect 161492 354 161520 818
rect 161266 326 161520 354
rect 160560 264 160612 270
rect 160560 206 160612 212
rect 161266 -960 161378 326
rect 161676 66 161704 2774
rect 163884 610 163912 2774
rect 164884 808 164936 814
rect 164884 750 164936 756
rect 163872 604 163924 610
rect 163872 546 163924 552
rect 164896 480 164924 750
rect 162308 264 162360 270
rect 162462 218 162574 480
rect 162360 212 162574 218
rect 162308 206 162574 212
rect 162320 190 162574 206
rect 161664 60 161716 66
rect 161664 2 161716 8
rect 162462 -960 162574 190
rect 163658 218 163770 480
rect 163658 202 163912 218
rect 163658 196 163924 202
rect 163658 190 163872 196
rect 163658 -960 163770 190
rect 163872 138 163924 144
rect 164854 -960 164966 480
rect 165080 406 165108 2774
rect 165908 2774 166166 2802
rect 165908 474 165936 2774
rect 166172 740 166224 746
rect 166172 682 166224 688
rect 166184 626 166212 682
rect 167012 678 167040 2858
rect 167242 2802 167270 3060
rect 168346 2802 168374 3060
rect 169450 2922 169478 3060
rect 170554 2922 170582 3060
rect 169438 2916 169490 2922
rect 169438 2858 169490 2864
rect 169576 2916 169628 2922
rect 169576 2858 169628 2864
rect 170542 2916 170594 2922
rect 170542 2858 170594 2864
rect 167242 2774 167408 2802
rect 166092 598 166212 626
rect 167000 672 167052 678
rect 167000 614 167052 620
rect 167184 672 167236 678
rect 167184 614 167236 620
rect 166092 480 166120 598
rect 167196 480 167224 614
rect 165896 468 165948 474
rect 165896 410 165948 416
rect 165068 400 165120 406
rect 165068 342 165120 348
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 167380 134 167408 2774
rect 168208 2774 168374 2802
rect 168208 338 168236 2774
rect 169588 882 169616 2858
rect 171658 2802 171686 3060
rect 172762 2802 172790 3060
rect 172980 2916 173032 2922
rect 172980 2858 173032 2864
rect 171612 2774 171686 2802
rect 172716 2774 172790 2802
rect 169576 876 169628 882
rect 169576 818 169628 824
rect 169576 672 169628 678
rect 168392 598 168604 626
rect 169576 614 169628 620
rect 168392 480 168420 598
rect 168196 332 168248 338
rect 168196 274 168248 280
rect 167368 128 167420 134
rect 167368 70 167420 76
rect 168350 -960 168462 480
rect 168576 354 168604 598
rect 169588 480 169616 614
rect 168576 326 168696 354
rect 168668 134 168696 326
rect 168656 128 168708 134
rect 168656 70 168708 76
rect 169546 -960 169658 480
rect 170588 400 170640 406
rect 170742 354 170854 480
rect 170640 348 170854 354
rect 170588 342 170854 348
rect 170600 326 170854 342
rect 170742 -960 170854 326
rect 171612 270 171640 2774
rect 171938 354 172050 480
rect 172152 468 172204 474
rect 172152 410 172204 416
rect 172164 354 172192 410
rect 171938 326 172192 354
rect 171600 264 171652 270
rect 171600 206 171652 212
rect 171938 -960 172050 326
rect 172716 202 172744 2774
rect 172992 746 173020 2858
rect 173866 2802 173894 3060
rect 174970 2922 174998 3060
rect 174958 2916 175010 2922
rect 174958 2858 175010 2864
rect 175280 2916 175332 2922
rect 175280 2858 175332 2864
rect 173820 2774 173894 2802
rect 173820 814 173848 2774
rect 173808 808 173860 814
rect 173808 750 173860 756
rect 172980 740 173032 746
rect 172980 682 173032 688
rect 173164 740 173216 746
rect 173164 682 173216 688
rect 173176 480 173204 682
rect 175292 678 175320 2858
rect 176074 2802 176102 3060
rect 177178 2802 177206 3060
rect 178282 2922 178310 3060
rect 178270 2916 178322 2922
rect 178270 2858 178322 2864
rect 179386 2802 179414 3060
rect 179512 2916 179564 2922
rect 179512 2858 179564 2864
rect 176028 2774 176102 2802
rect 177132 2774 177206 2802
rect 179340 2774 179414 2802
rect 175280 672 175332 678
rect 175280 614 175332 620
rect 174268 604 174320 610
rect 174268 546 174320 552
rect 174280 480 174308 546
rect 172704 196 172756 202
rect 172704 138 172756 144
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 218 175546 480
rect 176028 338 176056 2774
rect 176660 604 176712 610
rect 176660 546 176712 552
rect 176672 480 176700 546
rect 176016 332 176068 338
rect 176016 274 176068 280
rect 175434 202 175688 218
rect 175434 196 175700 202
rect 175434 190 175648 196
rect 175434 -960 175546 190
rect 175648 138 175700 144
rect 176630 -960 176742 480
rect 177132 134 177160 2774
rect 178040 536 178092 542
rect 177826 354 177938 480
rect 178040 478 178092 484
rect 178052 354 178080 478
rect 179022 354 179134 480
rect 179340 406 179368 2774
rect 179524 746 179552 2858
rect 180490 2802 180518 3060
rect 181594 2922 181622 3060
rect 182698 2922 182726 3060
rect 181582 2916 181634 2922
rect 181582 2858 181634 2864
rect 181720 2916 181772 2922
rect 181720 2858 181772 2864
rect 182686 2916 182738 2922
rect 182686 2858 182738 2864
rect 180444 2774 180518 2802
rect 179512 740 179564 746
rect 179512 682 179564 688
rect 177826 326 178080 354
rect 178880 338 179134 354
rect 179328 400 179380 406
rect 179328 342 179380 348
rect 178868 332 179134 338
rect 177120 128 177172 134
rect 177120 70 177172 76
rect 177826 -960 177938 326
rect 178920 326 179134 332
rect 178868 274 178920 280
rect 179022 -960 179134 326
rect 180218 82 180330 480
rect 180444 474 180472 2774
rect 181444 740 181496 746
rect 181444 682 181496 688
rect 181456 480 181484 682
rect 181732 678 181760 2858
rect 183802 2802 183830 3060
rect 184906 2802 184934 3060
rect 186010 2802 186038 3060
rect 187114 2802 187142 3060
rect 187700 2916 187752 2922
rect 187700 2858 187752 2864
rect 183572 2774 183830 2802
rect 184860 2774 184934 2802
rect 185964 2774 186038 2802
rect 187068 2774 187142 2802
rect 181720 672 181772 678
rect 181720 614 181772 620
rect 182548 672 182600 678
rect 182548 614 182600 620
rect 182560 480 182588 614
rect 180432 468 180484 474
rect 180432 410 180484 416
rect 180432 128 180484 134
rect 180218 76 180432 82
rect 180218 70 180484 76
rect 180218 54 180472 70
rect 180218 -960 180330 54
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183572 202 183600 2774
rect 183744 876 183796 882
rect 183744 818 183796 824
rect 183756 480 183784 818
rect 184860 610 184888 2774
rect 184940 808 184992 814
rect 184940 750 184992 756
rect 184848 604 184900 610
rect 184848 546 184900 552
rect 184952 480 184980 750
rect 185964 542 185992 2774
rect 185952 536 186004 542
rect 183560 196 183612 202
rect 183560 138 183612 144
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 185952 478 186004 484
rect 186106 218 186218 480
rect 187068 338 187096 2774
rect 187712 746 187740 2858
rect 188218 2802 188246 3060
rect 189322 2922 189350 3060
rect 189310 2916 189362 2922
rect 189310 2858 189362 2864
rect 190426 2802 190454 3060
rect 191530 2802 191558 3060
rect 192634 2802 192662 3060
rect 193738 2802 193766 3060
rect 194842 2802 194870 3060
rect 195946 2802 195974 3060
rect 197050 2802 197078 3060
rect 198154 2802 198182 3060
rect 188172 2774 188246 2802
rect 190380 2774 190454 2802
rect 191484 2774 191558 2802
rect 192588 2774 192662 2802
rect 193692 2774 193766 2802
rect 194796 2774 194870 2802
rect 195900 2774 195974 2802
rect 197004 2774 197078 2802
rect 198108 2774 198182 2802
rect 199258 2802 199286 3060
rect 200362 2802 200390 3060
rect 201466 2802 201494 3060
rect 202570 2802 202598 3060
rect 203674 2802 203702 3060
rect 199258 2774 199332 2802
rect 187700 740 187752 746
rect 187700 682 187752 688
rect 187056 332 187108 338
rect 187056 274 187108 280
rect 186320 264 186372 270
rect 186106 212 186320 218
rect 187302 218 187414 480
rect 186106 206 186372 212
rect 186106 190 186360 206
rect 187160 202 187414 218
rect 187148 196 187414 202
rect 186106 -960 186218 190
rect 187200 190 187414 196
rect 187148 138 187200 144
rect 187302 -960 187414 190
rect 188172 134 188200 2774
rect 190380 746 190408 2774
rect 190828 944 190880 950
rect 190828 886 190880 892
rect 190368 740 190420 746
rect 190368 682 190420 688
rect 188528 672 188580 678
rect 188528 614 188580 620
rect 188540 480 188568 614
rect 189724 604 189776 610
rect 189724 546 189776 552
rect 189736 480 189764 546
rect 190840 480 190868 886
rect 191484 882 191512 2774
rect 191472 876 191524 882
rect 191472 818 191524 824
rect 192588 814 192616 2774
rect 192576 808 192628 814
rect 192576 750 192628 756
rect 193220 808 193272 814
rect 193220 750 193272 756
rect 193232 480 193260 750
rect 188160 128 188212 134
rect 188160 70 188212 76
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 354 192106 480
rect 192208 468 192260 474
rect 192208 410 192260 416
rect 192220 354 192248 410
rect 191994 326 192248 354
rect 191994 -960 192106 326
rect 193190 -960 193302 480
rect 193692 270 193720 2774
rect 194416 740 194468 746
rect 194416 682 194468 688
rect 194428 480 194456 682
rect 193680 264 193732 270
rect 193680 206 193732 212
rect 194386 -960 194498 480
rect 194796 202 194824 2774
rect 195612 672 195664 678
rect 195612 614 195664 620
rect 195624 480 195652 614
rect 195900 610 195928 2774
rect 195888 604 195940 610
rect 195888 546 195940 552
rect 197004 542 197032 2774
rect 198108 950 198136 2774
rect 198096 944 198148 950
rect 198096 886 198148 892
rect 196992 536 197044 542
rect 194784 196 194836 202
rect 194784 138 194836 144
rect 195582 -960 195694 480
rect 196778 354 196890 480
rect 196992 478 197044 484
rect 196992 400 197044 406
rect 196778 348 196992 354
rect 196778 342 197044 348
rect 196778 326 197032 342
rect 196778 -960 196890 326
rect 197882 218 197994 480
rect 198096 264 198148 270
rect 197882 212 198096 218
rect 199078 218 199190 480
rect 199304 474 199332 2774
rect 200316 2774 200390 2802
rect 201420 2774 201494 2802
rect 202524 2774 202598 2802
rect 203628 2774 203702 2802
rect 204260 2848 204312 2854
rect 204778 2802 204806 3060
rect 205640 2916 205692 2922
rect 205640 2858 205692 2864
rect 204260 2790 204312 2796
rect 200316 814 200344 2774
rect 200304 808 200356 814
rect 200304 750 200356 756
rect 201420 746 201448 2774
rect 201408 740 201460 746
rect 201408 682 201460 688
rect 201500 740 201552 746
rect 201500 682 201552 688
rect 200304 604 200356 610
rect 200304 546 200356 552
rect 200316 480 200344 546
rect 201512 480 201540 682
rect 202524 678 202552 2774
rect 202512 672 202564 678
rect 202512 614 202564 620
rect 202696 604 202748 610
rect 202696 546 202748 552
rect 202708 480 202736 546
rect 199292 468 199344 474
rect 199292 410 199344 416
rect 197882 206 198148 212
rect 197882 190 198136 206
rect 198936 202 199190 218
rect 198924 196 199190 202
rect 197882 -960 197994 190
rect 198976 190 199190 196
rect 198924 138 198976 144
rect 199078 -960 199190 190
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203628 406 203656 2774
rect 203892 808 203944 814
rect 203892 750 203944 756
rect 203904 480 203932 750
rect 204272 678 204300 2790
rect 204732 2774 204806 2802
rect 204260 672 204312 678
rect 204260 614 204312 620
rect 203616 400 203668 406
rect 203616 342 203668 348
rect 203862 -960 203974 480
rect 204732 270 204760 2774
rect 205652 746 205680 2858
rect 205882 2802 205910 3060
rect 206986 2854 207014 3060
rect 208090 2922 208118 3060
rect 208078 2916 208130 2922
rect 208078 2858 208130 2864
rect 205836 2774 205910 2802
rect 206974 2848 207026 2854
rect 209194 2802 209222 3060
rect 210298 2802 210326 3060
rect 211402 2802 211430 3060
rect 211620 2916 211672 2922
rect 211620 2858 211672 2864
rect 206974 2790 207026 2796
rect 209148 2774 209222 2802
rect 210252 2774 210326 2802
rect 211356 2774 211430 2802
rect 205640 740 205692 746
rect 205640 682 205692 688
rect 205058 354 205170 480
rect 205058 338 205312 354
rect 205058 332 205324 338
rect 205058 326 205272 332
rect 204720 264 204772 270
rect 204720 206 204772 212
rect 205058 -960 205170 326
rect 205272 274 205324 280
rect 205836 202 205864 2774
rect 207388 672 207440 678
rect 207388 614 207440 620
rect 207400 480 207428 614
rect 209148 610 209176 2774
rect 210252 814 210280 2774
rect 210976 876 211028 882
rect 210976 818 211028 824
rect 210240 808 210292 814
rect 210240 750 210292 756
rect 209780 740 209832 746
rect 209780 682 209832 688
rect 209136 604 209188 610
rect 209136 546 209188 552
rect 209792 480 209820 682
rect 210988 480 211016 818
rect 206162 218 206274 480
rect 206376 264 206428 270
rect 206162 212 206376 218
rect 206162 206 206428 212
rect 205824 196 205876 202
rect 205824 138 205876 144
rect 206162 190 206416 206
rect 206162 -960 206274 190
rect 207358 -960 207470 480
rect 208554 354 208666 480
rect 208768 400 208820 406
rect 208554 348 208768 354
rect 208554 342 208820 348
rect 208554 326 208808 342
rect 208554 -960 208666 326
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211356 338 211384 2774
rect 211632 678 211660 2858
rect 212506 2802 212534 3060
rect 213610 2922 213638 3060
rect 214714 2922 214742 3060
rect 215818 2922 215846 3060
rect 213598 2916 213650 2922
rect 213598 2858 213650 2864
rect 213736 2916 213788 2922
rect 213736 2858 213788 2864
rect 214702 2916 214754 2922
rect 214702 2858 214754 2864
rect 214840 2916 214892 2922
rect 214840 2858 214892 2864
rect 215806 2916 215858 2922
rect 215806 2858 215858 2864
rect 216680 2916 216732 2922
rect 216680 2858 216732 2864
rect 212460 2774 212534 2802
rect 211620 672 211672 678
rect 211620 614 211672 620
rect 212172 672 212224 678
rect 212172 614 212224 620
rect 212184 480 212212 614
rect 211344 332 211396 338
rect 211344 274 211396 280
rect 212142 -960 212254 480
rect 212460 270 212488 2774
rect 213368 604 213420 610
rect 213368 546 213420 552
rect 213380 480 213408 546
rect 212448 264 212500 270
rect 212448 206 212500 212
rect 213338 -960 213450 480
rect 213748 406 213776 2858
rect 214472 808 214524 814
rect 214472 750 214524 756
rect 214484 480 214512 750
rect 214852 746 214880 2858
rect 215300 2848 215352 2854
rect 215300 2790 215352 2796
rect 214840 740 214892 746
rect 214840 682 214892 688
rect 215312 678 215340 2790
rect 215668 740 215720 746
rect 215668 682 215720 688
rect 215300 672 215352 678
rect 215300 614 215352 620
rect 215680 480 215708 682
rect 216692 610 216720 2858
rect 216922 2802 216950 3060
rect 218026 2938 218054 3060
rect 217980 2910 218054 2938
rect 219130 2922 219158 3060
rect 219118 2916 219170 2922
rect 217980 2854 218008 2910
rect 219118 2858 219170 2864
rect 220234 2854 220262 3060
rect 221338 2922 221366 3060
rect 222442 2922 222470 3060
rect 220360 2916 220412 2922
rect 220360 2858 220412 2864
rect 221326 2916 221378 2922
rect 221326 2858 221378 2864
rect 221464 2916 221516 2922
rect 221464 2858 221516 2864
rect 222430 2916 222482 2922
rect 222430 2858 222482 2864
rect 222568 2916 222620 2922
rect 222568 2858 222620 2864
rect 216876 2774 216950 2802
rect 217968 2848 218020 2854
rect 217968 2790 218020 2796
rect 218060 2848 218112 2854
rect 218060 2790 218112 2796
rect 220222 2848 220274 2854
rect 220222 2790 220274 2796
rect 216876 882 216904 2774
rect 216864 876 216916 882
rect 216864 818 216916 824
rect 218072 814 218100 2790
rect 218060 808 218112 814
rect 218060 750 218112 756
rect 220372 746 220400 2858
rect 220360 740 220412 746
rect 220360 682 220412 688
rect 220452 740 220504 746
rect 220452 682 220504 688
rect 216864 672 216916 678
rect 216864 614 216916 620
rect 216680 604 216732 610
rect 216680 546 216732 552
rect 216876 480 216904 614
rect 218060 604 218112 610
rect 218060 546 218112 552
rect 218072 480 218100 546
rect 220464 480 220492 682
rect 221476 678 221504 2858
rect 221464 672 221516 678
rect 221464 614 221516 620
rect 221556 604 221608 610
rect 221556 546 221608 552
rect 221568 480 221596 546
rect 213736 400 213788 406
rect 213736 342 213788 348
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 354 219338 480
rect 219440 400 219492 406
rect 219226 348 219440 354
rect 219226 342 219492 348
rect 219226 326 219480 342
rect 219226 -960 219338 326
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222580 406 222608 2858
rect 223546 2802 223574 3060
rect 224650 2922 224678 3060
rect 225754 2922 225782 3060
rect 224638 2916 224690 2922
rect 224638 2858 224690 2864
rect 224776 2916 224828 2922
rect 224776 2858 224828 2864
rect 225742 2916 225794 2922
rect 225742 2858 225794 2864
rect 226524 2916 226576 2922
rect 226524 2858 226576 2864
rect 223500 2774 223574 2802
rect 222568 400 222620 406
rect 222568 342 222620 348
rect 222722 354 222834 480
rect 222936 400 222988 406
rect 222722 348 222936 354
rect 222722 342 222988 348
rect 222722 326 222976 342
rect 222722 -960 222834 326
rect 223500 202 223528 2774
rect 223948 808 224000 814
rect 223948 750 224000 756
rect 223960 480 223988 750
rect 224788 746 224816 2858
rect 224960 2848 225012 2854
rect 224960 2790 225012 2796
rect 224776 740 224828 746
rect 224776 682 224828 688
rect 224972 610 225000 2790
rect 226340 672 226392 678
rect 226340 614 226392 620
rect 224960 604 225012 610
rect 224960 546 225012 552
rect 226352 480 226380 614
rect 223488 196 223540 202
rect 223488 138 223540 144
rect 223918 -960 224030 480
rect 225114 354 225226 480
rect 225328 468 225380 474
rect 225328 410 225380 416
rect 225340 354 225368 410
rect 225114 326 225368 354
rect 225114 -960 225226 326
rect 226310 -960 226422 480
rect 226536 406 226564 2858
rect 226858 2854 226886 3060
rect 227962 2922 227990 3060
rect 227950 2916 228002 2922
rect 227950 2858 228002 2864
rect 226846 2848 226898 2854
rect 229066 2802 229094 3060
rect 230170 2802 230198 3060
rect 230572 2916 230624 2922
rect 230572 2858 230624 2864
rect 226846 2790 226898 2796
rect 229020 2774 229094 2802
rect 230124 2774 230198 2802
rect 229020 814 229048 2774
rect 229008 808 229060 814
rect 229008 750 229060 756
rect 229836 808 229888 814
rect 229836 750 229888 756
rect 227536 604 227588 610
rect 227536 546 227588 552
rect 227548 480 227576 546
rect 229848 480 229876 750
rect 226524 400 226576 406
rect 226524 342 226576 348
rect 227506 -960 227618 480
rect 228548 128 228600 134
rect 228702 82 228814 480
rect 228600 76 228814 82
rect 228548 70 228814 76
rect 228560 54 228814 70
rect 228702 -960 228814 54
rect 229806 -960 229918 480
rect 230124 474 230152 2774
rect 230584 610 230612 2858
rect 231274 2802 231302 3060
rect 232378 2922 232406 3060
rect 233482 2922 233510 3060
rect 232366 2916 232418 2922
rect 232366 2858 232418 2864
rect 232504 2916 232556 2922
rect 232504 2858 232556 2864
rect 233470 2916 233522 2922
rect 233470 2858 233522 2864
rect 231228 2774 231302 2802
rect 231228 678 231256 2774
rect 231216 672 231268 678
rect 231216 614 231268 620
rect 230572 604 230624 610
rect 230572 546 230624 552
rect 232228 604 232280 610
rect 232228 546 232280 552
rect 232240 480 232268 546
rect 230112 468 230164 474
rect 230112 410 230164 416
rect 231002 354 231114 480
rect 231216 400 231268 406
rect 231002 348 231216 354
rect 231002 342 231268 348
rect 231002 326 231256 342
rect 231002 -960 231114 326
rect 232198 -960 232310 480
rect 232516 134 232544 2858
rect 234586 2802 234614 3060
rect 234712 2916 234764 2922
rect 234712 2858 234764 2864
rect 234540 2774 234614 2802
rect 234540 814 234568 2774
rect 234528 808 234580 814
rect 234528 750 234580 756
rect 233424 740 233476 746
rect 233424 682 233476 688
rect 233436 480 233464 682
rect 234620 672 234672 678
rect 234620 614 234672 620
rect 234632 480 234660 614
rect 234724 610 234752 2858
rect 235690 2802 235718 3060
rect 236794 2922 236822 3060
rect 236782 2916 236834 2922
rect 236782 2858 236834 2864
rect 237898 2802 237926 3060
rect 239002 2802 239030 3060
rect 240106 2802 240134 3060
rect 241210 2802 241238 3060
rect 242314 2802 242342 3060
rect 242900 2916 242952 2922
rect 242900 2858 242952 2864
rect 235644 2774 235718 2802
rect 237852 2774 237926 2802
rect 238956 2774 239030 2802
rect 240060 2774 240134 2802
rect 241164 2774 241238 2802
rect 242268 2774 242342 2802
rect 234712 604 234764 610
rect 234712 546 234764 552
rect 232504 128 232556 134
rect 232504 70 232556 76
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235644 406 235672 2774
rect 237852 746 237880 2774
rect 237840 740 237892 746
rect 237840 682 237892 688
rect 238956 678 238984 2774
rect 238944 672 238996 678
rect 238944 614 238996 620
rect 237012 604 237064 610
rect 237012 546 237064 552
rect 237024 480 237052 546
rect 235632 400 235684 406
rect 235632 342 235684 348
rect 235786 354 235898 480
rect 236000 400 236052 406
rect 235786 348 236000 354
rect 235786 342 236052 348
rect 235786 326 236040 342
rect 235786 -960 235898 326
rect 236982 -960 237094 480
rect 237932 264 237984 270
rect 238086 218 238198 480
rect 237984 212 238198 218
rect 237932 206 238198 212
rect 237944 190 238198 206
rect 238086 -960 238198 190
rect 239282 354 239394 480
rect 239496 468 239548 474
rect 239496 410 239548 416
rect 239508 354 239536 410
rect 240060 406 240088 2774
rect 240508 672 240560 678
rect 240508 614 240560 620
rect 240520 480 240548 614
rect 241164 610 241192 2774
rect 241152 604 241204 610
rect 241152 546 241204 552
rect 241704 604 241756 610
rect 241704 546 241756 552
rect 241716 480 241744 546
rect 239282 326 239536 354
rect 240048 400 240100 406
rect 240048 342 240100 348
rect 239282 -960 239394 326
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242268 270 242296 2774
rect 242912 480 242940 2858
rect 243418 2802 243446 3060
rect 244522 2802 244550 3060
rect 245626 2802 245654 3060
rect 246730 2922 246758 3060
rect 246718 2916 246770 2922
rect 246718 2858 246770 2864
rect 247592 2916 247644 2922
rect 247592 2858 247644 2864
rect 243372 2774 243446 2802
rect 244476 2774 244550 2802
rect 245580 2774 245654 2802
rect 242256 264 242308 270
rect 242256 206 242308 212
rect 242870 -960 242982 480
rect 243372 474 243400 2774
rect 244476 678 244504 2774
rect 244464 672 244516 678
rect 244464 614 244516 620
rect 245200 672 245252 678
rect 245200 614 245252 620
rect 245212 480 245240 614
rect 245580 610 245608 2774
rect 245568 604 245620 610
rect 245568 546 245620 552
rect 246396 604 246448 610
rect 246396 546 246448 552
rect 246408 480 246436 546
rect 247604 480 247632 2858
rect 247834 2802 247862 3060
rect 248938 2802 248966 3060
rect 247788 2774 247862 2802
rect 248892 2774 248966 2802
rect 249892 2848 249944 2854
rect 249892 2790 249944 2796
rect 250042 2802 250070 3060
rect 251146 2922 251174 3060
rect 251134 2916 251186 2922
rect 251134 2858 251186 2864
rect 252250 2802 252278 3060
rect 253354 2854 253382 3060
rect 253480 2916 253532 2922
rect 253480 2858 253532 2864
rect 243360 468 243412 474
rect 243360 410 243412 416
rect 244066 354 244178 480
rect 244280 400 244332 406
rect 244066 348 244280 354
rect 244066 342 244332 348
rect 244066 326 244320 342
rect 244066 -960 244178 326
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 247788 406 247816 2774
rect 248788 740 248840 746
rect 248788 682 248840 688
rect 248800 480 248828 682
rect 248892 678 248920 2774
rect 248880 672 248932 678
rect 248880 614 248932 620
rect 249904 626 249932 2790
rect 250042 2774 250116 2802
rect 249904 598 250024 626
rect 250088 610 250116 2774
rect 252204 2774 252278 2802
rect 253342 2848 253394 2854
rect 253342 2790 253394 2796
rect 252204 746 252232 2774
rect 252192 740 252244 746
rect 252192 682 252244 688
rect 249996 480 250024 598
rect 250076 604 250128 610
rect 250076 546 250128 552
rect 251180 604 251232 610
rect 251180 546 251232 552
rect 251192 480 251220 546
rect 253492 480 253520 2858
rect 254458 2802 254486 3060
rect 255562 2802 255590 3060
rect 256666 2922 256694 3060
rect 256654 2916 256706 2922
rect 256654 2858 256706 2864
rect 257068 2916 257120 2922
rect 257068 2858 257120 2864
rect 254412 2774 254486 2802
rect 255516 2774 255590 2802
rect 254412 610 254440 2774
rect 254400 604 254452 610
rect 254400 546 254452 552
rect 254676 604 254728 610
rect 254676 546 254728 552
rect 254688 480 254716 546
rect 247776 400 247828 406
rect 247776 342 247828 348
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 354 252458 480
rect 252560 400 252612 406
rect 252346 348 252560 354
rect 252346 342 252612 348
rect 252346 326 252600 342
rect 252346 -960 252458 326
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255516 406 255544 2774
rect 257080 480 257108 2858
rect 257770 2802 257798 3060
rect 258874 2802 258902 3060
rect 259978 2922 260006 3060
rect 259966 2916 260018 2922
rect 259966 2858 260018 2864
rect 257724 2774 257798 2802
rect 258828 2774 258902 2802
rect 259460 2848 259512 2854
rect 261082 2802 261110 3060
rect 261760 2916 261812 2922
rect 261760 2858 261812 2864
rect 259460 2790 259512 2796
rect 257724 610 257752 2774
rect 257712 604 257764 610
rect 257712 546 257764 552
rect 258264 604 258316 610
rect 258264 546 258316 552
rect 258276 480 258304 546
rect 255504 400 255556 406
rect 255504 342 255556 348
rect 255842 354 255954 480
rect 256056 400 256108 406
rect 255842 348 256056 354
rect 255842 342 256108 348
rect 255842 326 256096 342
rect 255842 -960 255954 326
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 258828 406 258856 2774
rect 259472 480 259500 2790
rect 261036 2774 261110 2802
rect 261036 610 261064 2774
rect 261024 604 261076 610
rect 261024 546 261076 552
rect 261772 480 261800 2858
rect 262186 2854 262214 3060
rect 262174 2848 262226 2854
rect 263290 2802 263318 3060
rect 264394 2922 264422 3060
rect 264382 2916 264434 2922
rect 264382 2858 264434 2864
rect 265348 2916 265400 2922
rect 265348 2858 265400 2864
rect 262174 2790 262226 2796
rect 263244 2774 263318 2802
rect 262956 672 263008 678
rect 262956 614 263008 620
rect 262968 480 262996 614
rect 258816 400 258868 406
rect 258816 342 258868 348
rect 259430 -960 259542 480
rect 260626 354 260738 480
rect 260840 400 260892 406
rect 260626 348 260840 354
rect 260626 342 260892 348
rect 260626 326 260880 342
rect 260626 -960 260738 326
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 263244 406 263272 2774
rect 264152 604 264204 610
rect 264152 546 264204 552
rect 264164 480 264192 546
rect 265360 480 265388 2858
rect 265498 2802 265526 3060
rect 266602 2938 266630 3060
rect 266602 2910 266676 2938
rect 267706 2922 267734 3060
rect 265452 2774 265526 2802
rect 266544 2848 266596 2854
rect 266544 2790 266596 2796
rect 265452 678 265480 2774
rect 265440 672 265492 678
rect 265440 614 265492 620
rect 266556 480 266584 2790
rect 266648 610 266676 2910
rect 267694 2916 267746 2922
rect 267694 2858 267746 2864
rect 267832 2916 267884 2922
rect 267832 2858 267884 2864
rect 267844 1578 267872 2858
rect 268810 2854 268838 3060
rect 269914 2922 269942 3060
rect 269902 2916 269954 2922
rect 269902 2858 269954 2864
rect 268798 2848 268850 2854
rect 271018 2802 271046 3060
rect 271236 2916 271288 2922
rect 271236 2858 271288 2864
rect 268798 2790 268850 2796
rect 267752 1550 267872 1578
rect 270972 2774 271046 2802
rect 266636 604 266688 610
rect 266636 546 266688 552
rect 267752 480 267780 1550
rect 270972 610 271000 2774
rect 268844 604 268896 610
rect 268844 546 268896 552
rect 270960 604 271012 610
rect 270960 546 271012 552
rect 268856 480 268884 546
rect 271248 480 271276 2858
rect 272122 2802 272150 3060
rect 273226 2922 273254 3060
rect 273214 2916 273266 2922
rect 273214 2858 273266 2864
rect 273628 2916 273680 2922
rect 273628 2858 273680 2864
rect 272076 2774 272150 2802
rect 272432 2848 272484 2854
rect 272432 2790 272484 2796
rect 263232 400 263284 406
rect 263232 342 263284 348
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 354 270122 480
rect 270224 400 270276 406
rect 270010 348 270224 354
rect 270010 342 270276 348
rect 270010 326 270264 342
rect 270010 -960 270122 326
rect 271206 -960 271318 480
rect 272076 406 272104 2774
rect 272444 480 272472 2790
rect 273640 480 273668 2858
rect 274330 2854 274358 3060
rect 275434 2922 275462 3060
rect 275422 2916 275474 2922
rect 275422 2858 275474 2864
rect 276020 2916 276072 2922
rect 276020 2858 276072 2864
rect 274318 2848 274370 2854
rect 274318 2790 274370 2796
rect 274824 2848 274876 2854
rect 274824 2790 274876 2796
rect 274836 480 274864 2790
rect 276032 480 276060 2858
rect 276538 2854 276566 3060
rect 277642 2922 277670 3060
rect 277630 2916 277682 2922
rect 277630 2858 277682 2864
rect 278320 2916 278372 2922
rect 278320 2858 278372 2864
rect 276526 2848 276578 2854
rect 276526 2790 276578 2796
rect 277124 604 277176 610
rect 277124 546 277176 552
rect 277136 480 277164 546
rect 278332 480 278360 2858
rect 278746 2802 278774 3060
rect 279850 2922 279878 3060
rect 279838 2916 279890 2922
rect 279838 2858 279890 2864
rect 280712 2916 280764 2922
rect 280712 2858 280764 2864
rect 278700 2774 278774 2802
rect 279516 2848 279568 2854
rect 279516 2790 279568 2796
rect 278700 610 278728 2774
rect 278688 604 278740 610
rect 278688 546 278740 552
rect 279528 480 279556 2790
rect 280724 480 280752 2858
rect 280954 2854 280982 3060
rect 282058 2922 282086 3060
rect 283162 2922 283190 3060
rect 282046 2916 282098 2922
rect 282046 2858 282098 2864
rect 283150 2916 283202 2922
rect 283150 2858 283202 2864
rect 280942 2848 280994 2854
rect 280942 2790 280994 2796
rect 281908 2848 281960 2854
rect 284266 2802 284294 3060
rect 285370 2938 285398 3060
rect 281908 2790 281960 2796
rect 281920 480 281948 2790
rect 283300 2774 284294 2802
rect 284404 2910 285398 2938
rect 283300 1578 283328 2774
rect 284404 1578 284432 2910
rect 286474 2854 286502 3060
rect 287578 2922 287606 3060
rect 288682 2922 288710 3060
rect 286600 2916 286652 2922
rect 286600 2858 286652 2864
rect 287566 2916 287618 2922
rect 287566 2858 287618 2864
rect 287796 2916 287848 2922
rect 287796 2858 287848 2864
rect 288670 2916 288722 2922
rect 288670 2858 288722 2864
rect 285404 2848 285456 2854
rect 285404 2790 285456 2796
rect 286462 2848 286514 2854
rect 286462 2790 286514 2796
rect 283116 1550 283328 1578
rect 284312 1550 284432 1578
rect 283116 480 283144 1550
rect 284312 480 284340 1550
rect 285416 480 285444 2790
rect 286612 480 286640 2858
rect 287808 480 287836 2858
rect 289786 2802 289814 3060
rect 290890 2802 290918 3060
rect 291994 2802 292022 3060
rect 293098 2802 293126 3060
rect 294202 2922 294230 3060
rect 293684 2916 293736 2922
rect 293684 2858 293736 2864
rect 294190 2916 294242 2922
rect 294190 2858 294242 2864
rect 289464 2774 289814 2802
rect 290200 2774 290918 2802
rect 291856 2774 292022 2802
rect 292592 2774 293126 2802
rect 272064 400 272116 406
rect 272064 342 272116 348
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 354 289074 480
rect 289464 354 289492 2774
rect 290200 480 290228 2774
rect 288962 326 289492 354
rect 288962 -960 289074 326
rect 290158 -960 290270 480
rect 291354 354 291466 480
rect 291856 354 291884 2774
rect 292592 480 292620 2774
rect 293696 480 293724 2858
rect 295306 2802 295334 3060
rect 296410 2802 296438 3060
rect 297514 2802 297542 3060
rect 298618 2802 298646 3060
rect 299722 2802 299750 3060
rect 300826 2802 300854 3060
rect 295260 2774 295334 2802
rect 296088 2774 296438 2802
rect 297468 2774 297542 2802
rect 298480 2774 298646 2802
rect 299676 2774 299750 2802
rect 300780 2774 300854 2802
rect 301930 2802 301958 3060
rect 303034 2802 303062 3060
rect 304138 2802 304166 3060
rect 305242 2802 305270 3060
rect 306346 2802 306374 3060
rect 301930 2774 302004 2802
rect 303034 2774 303200 2802
rect 304138 2774 304212 2802
rect 305242 2774 305592 2802
rect 291354 326 291884 354
rect 291354 -960 291466 326
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 354 294962 480
rect 295260 354 295288 2774
rect 296088 480 296116 2774
rect 294850 326 295288 354
rect 294850 -960 294962 326
rect 296046 -960 296158 480
rect 297242 354 297354 480
rect 297468 354 297496 2774
rect 298480 480 298508 2774
rect 299676 480 299704 2774
rect 300780 480 300808 2774
rect 301976 480 302004 2774
rect 303172 480 303200 2774
rect 297242 326 297496 354
rect 297242 -960 297354 326
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304184 354 304212 2774
rect 305564 480 305592 2774
rect 306300 2774 306374 2802
rect 307450 2802 307478 3060
rect 308554 2802 308582 3060
rect 309658 2802 309686 3060
rect 310762 2802 310790 3060
rect 311866 2802 311894 3060
rect 307450 2774 307524 2802
rect 308554 2774 309088 2802
rect 309658 2774 309824 2802
rect 310762 2774 311480 2802
rect 304326 354 304438 480
rect 304184 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306300 354 306328 2774
rect 307496 610 307524 2774
rect 307484 604 307536 610
rect 307484 546 307536 552
rect 307944 604 307996 610
rect 307944 546 307996 552
rect 307956 480 307984 546
rect 309060 480 309088 2774
rect 306718 354 306830 480
rect 306300 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 2774
rect 311452 480 311480 2774
rect 311820 2774 311894 2802
rect 312970 2802 312998 3060
rect 314074 2802 314102 3060
rect 315178 2802 315206 3060
rect 316282 2854 316310 3060
rect 317386 2938 317414 3060
rect 317248 2910 317414 2938
rect 316270 2848 316322 2854
rect 312970 2774 313044 2802
rect 314074 2774 314148 2802
rect 315178 2774 315252 2802
rect 316270 2790 316322 2796
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 311820 406 311848 2774
rect 313016 610 313044 2774
rect 313004 604 313056 610
rect 313004 546 313056 552
rect 313832 604 313884 610
rect 313832 546 313884 552
rect 313844 480 313872 546
rect 311808 400 311860 406
rect 311808 342 311860 348
rect 312452 400 312504 406
rect 312606 354 312718 480
rect 312504 348 312718 354
rect 312452 342 312718 348
rect 312464 326 312718 342
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314120 406 314148 2774
rect 315224 610 315252 2774
rect 317248 610 317276 2910
rect 317328 2848 317380 2854
rect 317328 2790 317380 2796
rect 318490 2802 318518 3060
rect 319594 2802 319622 3060
rect 320698 2922 320726 3060
rect 320686 2916 320738 2922
rect 320686 2858 320738 2864
rect 321802 2802 321830 3060
rect 322906 2922 322934 3060
rect 322112 2916 322164 2922
rect 322112 2858 322164 2864
rect 322894 2916 322946 2922
rect 322894 2858 322946 2864
rect 315212 604 315264 610
rect 315212 546 315264 552
rect 316224 604 316276 610
rect 316224 546 316276 552
rect 317236 604 317288 610
rect 317236 546 317288 552
rect 316236 480 316264 546
rect 317340 480 317368 2790
rect 318490 2774 318564 2802
rect 319594 2774 319668 2802
rect 321802 2774 321876 2802
rect 318536 746 318564 2774
rect 318524 740 318576 746
rect 318524 682 318576 688
rect 319640 610 319668 2774
rect 319720 740 319772 746
rect 319720 682 319772 688
rect 318524 604 318576 610
rect 318524 546 318576 552
rect 319628 604 319680 610
rect 319628 546 319680 552
rect 318536 480 318564 546
rect 319732 480 319760 682
rect 320916 604 320968 610
rect 320916 546 320968 552
rect 320928 480 320956 546
rect 314108 400 314160 406
rect 314108 342 314160 348
rect 314844 400 314896 406
rect 314998 354 315110 480
rect 314896 348 315110 354
rect 314844 342 315110 348
rect 314856 326 315110 342
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 321848 406 321876 2774
rect 322124 480 322152 2858
rect 324010 2802 324038 3060
rect 325114 2922 325142 3060
rect 324412 2916 324464 2922
rect 324412 2858 324464 2864
rect 325102 2916 325154 2922
rect 325102 2858 325154 2864
rect 324010 2774 324084 2802
rect 324056 610 324084 2774
rect 324044 604 324096 610
rect 324044 546 324096 552
rect 324424 480 324452 2858
rect 326218 2802 326246 3060
rect 326804 2916 326856 2922
rect 326804 2858 326856 2864
rect 326218 2774 326292 2802
rect 326264 610 326292 2774
rect 325608 604 325660 610
rect 325608 546 325660 552
rect 326252 604 326304 610
rect 326252 546 326304 552
rect 325620 480 325648 546
rect 326816 480 326844 2858
rect 327322 2802 327350 3060
rect 328426 2802 328454 3060
rect 329530 2922 329558 3060
rect 329518 2916 329570 2922
rect 329518 2858 329570 2864
rect 327322 2774 327396 2802
rect 321836 400 321888 406
rect 321836 342 321888 348
rect 322082 -960 322194 480
rect 323124 400 323176 406
rect 323278 354 323390 480
rect 323176 348 323390 354
rect 323124 342 323390 348
rect 323136 326 323390 342
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327368 406 327396 2774
rect 328380 2774 328454 2802
rect 330634 2802 330662 3060
rect 331738 2922 331766 3060
rect 331588 2916 331640 2922
rect 331588 2858 331640 2864
rect 331726 2916 331778 2922
rect 331726 2858 331778 2864
rect 330634 2774 330708 2802
rect 328380 610 328408 2774
rect 328000 604 328052 610
rect 328000 546 328052 552
rect 328368 604 328420 610
rect 328368 546 328420 552
rect 330392 604 330444 610
rect 330392 546 330444 552
rect 328012 480 328040 546
rect 330404 480 330432 546
rect 327356 400 327408 406
rect 327356 342 327408 348
rect 327970 -960 328082 480
rect 329012 400 329064 406
rect 329166 354 329278 480
rect 329064 348 329278 354
rect 329012 342 329278 348
rect 329024 326 329278 342
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 330680 406 330708 2774
rect 331600 480 331628 2858
rect 332842 2802 332870 3060
rect 333796 2916 333848 2922
rect 333796 2858 333848 2864
rect 332842 2774 332916 2802
rect 332888 610 332916 2774
rect 333808 1578 333836 2858
rect 333946 2802 333974 3060
rect 335050 2922 335078 3060
rect 335038 2916 335090 2922
rect 335038 2858 335090 2864
rect 336154 2854 336182 3060
rect 336464 2916 336516 2922
rect 336464 2858 336516 2864
rect 336142 2848 336194 2854
rect 333946 2774 334020 2802
rect 336142 2790 336194 2796
rect 333808 1550 333928 1578
rect 332876 604 332928 610
rect 332876 546 332928 552
rect 333900 480 333928 1550
rect 333992 678 334020 2774
rect 333980 672 334032 678
rect 333980 614 334032 620
rect 336280 672 336332 678
rect 336280 614 336332 620
rect 335084 604 335136 610
rect 335084 546 335136 552
rect 335096 480 335124 546
rect 336292 480 336320 614
rect 330668 400 330720 406
rect 330668 342 330720 348
rect 331558 -960 331670 480
rect 332508 400 332560 406
rect 332662 354 332774 480
rect 332560 348 332774 354
rect 332508 342 332774 348
rect 332520 326 332774 342
rect 332662 -960 332774 326
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 336476 406 336504 2858
rect 337258 2802 337286 3060
rect 338362 2802 338390 3060
rect 338672 2848 338724 2854
rect 337258 2774 337332 2802
rect 338362 2774 338436 2802
rect 338672 2790 338724 2796
rect 339466 2802 339494 3060
rect 340570 2922 340598 3060
rect 340558 2916 340610 2922
rect 340558 2858 340610 2864
rect 341674 2802 341702 3060
rect 342778 2854 342806 3060
rect 343364 2916 343416 2922
rect 343364 2858 343416 2864
rect 342766 2848 342818 2854
rect 337304 610 337332 2774
rect 337292 604 337344 610
rect 337292 546 337344 552
rect 336464 400 336516 406
rect 336464 342 336516 348
rect 337292 400 337344 406
rect 337446 354 337558 480
rect 338408 406 338436 2774
rect 338684 480 338712 2790
rect 339466 2774 339540 2802
rect 341674 2774 341748 2802
rect 342766 2790 342818 2796
rect 339512 678 339540 2774
rect 341720 746 341748 2774
rect 341708 740 341760 746
rect 341708 682 341760 688
rect 339500 672 339552 678
rect 339500 614 339552 620
rect 342168 672 342220 678
rect 342168 614 342220 620
rect 339868 604 339920 610
rect 339868 546 339920 552
rect 339880 480 339908 546
rect 342180 480 342208 614
rect 343376 480 343404 2858
rect 343882 2802 343910 3060
rect 344986 2904 345014 3060
rect 346090 2922 346118 3060
rect 346078 2916 346130 2922
rect 344986 2876 345060 2904
rect 345032 2802 345060 2876
rect 346078 2858 346130 2864
rect 347194 2854 347222 3060
rect 348298 2922 348326 3060
rect 347596 2916 347648 2922
rect 347596 2858 347648 2864
rect 348286 2916 348338 2922
rect 348286 2858 348338 2864
rect 343882 2774 343956 2802
rect 343928 610 343956 2774
rect 344940 2774 345060 2802
rect 345756 2848 345808 2854
rect 345756 2790 345808 2796
rect 347182 2848 347234 2854
rect 347182 2790 347234 2796
rect 344560 740 344612 746
rect 344560 682 344612 688
rect 343916 604 343968 610
rect 343916 546 343968 552
rect 344572 480 344600 682
rect 337344 348 337558 354
rect 337292 342 337558 348
rect 338396 400 338448 406
rect 338396 342 338448 348
rect 337304 326 337558 342
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340788 400 340840 406
rect 340942 354 341054 480
rect 340840 348 341054 354
rect 340788 342 341054 348
rect 340800 326 341054 342
rect 340942 -960 341054 326
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 344940 134 344968 2774
rect 345768 480 345796 2790
rect 346952 604 347004 610
rect 346952 546 347004 552
rect 346964 480 346992 546
rect 344928 128 344980 134
rect 344928 70 344980 76
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 347608 406 347636 2858
rect 349402 2854 349430 3060
rect 349896 2916 349948 2922
rect 349896 2858 349948 2864
rect 348792 2848 348844 2854
rect 348792 2790 348844 2796
rect 349390 2848 349442 2854
rect 349390 2790 349442 2796
rect 348804 610 348832 2790
rect 349908 678 349936 2858
rect 350506 2802 350534 3060
rect 350460 2774 350534 2802
rect 351610 2802 351638 3060
rect 352714 2922 352742 3060
rect 352702 2916 352754 2922
rect 352702 2858 352754 2864
rect 352840 2848 352892 2854
rect 351610 2774 351684 2802
rect 352840 2790 352892 2796
rect 353818 2802 353846 3060
rect 354922 2854 354950 3060
rect 356026 2938 356054 3060
rect 355784 2916 355836 2922
rect 355784 2858 355836 2864
rect 355888 2910 356054 2938
rect 354910 2848 354962 2854
rect 350460 746 350488 2774
rect 351656 814 351684 2774
rect 351644 808 351696 814
rect 351644 750 351696 756
rect 350448 740 350500 746
rect 350448 682 350500 688
rect 349896 672 349948 678
rect 349896 614 349948 620
rect 351644 672 351696 678
rect 351644 614 351696 620
rect 348792 604 348844 610
rect 348792 546 348844 552
rect 350448 604 350500 610
rect 350448 546 350500 552
rect 350460 480 350488 546
rect 351656 480 351684 614
rect 352852 480 352880 2790
rect 353818 2774 353892 2802
rect 354910 2790 354962 2796
rect 347596 400 347648 406
rect 347596 342 347648 348
rect 348026 82 348138 480
rect 349068 400 349120 406
rect 349222 354 349334 480
rect 349120 348 349334 354
rect 349068 342 349334 348
rect 349080 326 349334 342
rect 348240 128 348292 134
rect 348026 76 348240 82
rect 348026 70 348292 76
rect 348026 54 348280 70
rect 348026 -960 348138 54
rect 349222 -960 349334 326
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353864 270 353892 2774
rect 355232 808 355284 814
rect 355232 750 355284 756
rect 354036 740 354088 746
rect 354036 682 354088 688
rect 354048 480 354076 682
rect 355244 480 355272 750
rect 355796 610 355824 2858
rect 355784 604 355836 610
rect 355784 546 355836 552
rect 353852 264 353904 270
rect 353852 206 353904 212
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 355888 406 355916 2910
rect 357130 2802 357158 3060
rect 358234 2922 358262 3060
rect 358222 2916 358274 2922
rect 358222 2858 358274 2864
rect 359338 2854 359366 3060
rect 360108 2916 360160 2922
rect 360108 2858 360160 2864
rect 358728 2848 358780 2854
rect 357130 2774 357204 2802
rect 358728 2790 358780 2796
rect 359326 2848 359378 2854
rect 359326 2790 359378 2796
rect 357176 610 357204 2774
rect 356336 604 356388 610
rect 356336 546 356388 552
rect 357164 604 357216 610
rect 357164 546 357216 552
rect 356348 480 356376 546
rect 358740 480 358768 2790
rect 355876 400 355928 406
rect 355876 342 355928 348
rect 356306 -960 356418 480
rect 357348 264 357400 270
rect 357502 218 357614 480
rect 357400 212 357614 218
rect 357348 206 357614 212
rect 357360 190 357614 206
rect 357502 -960 357614 190
rect 358698 -960 358810 480
rect 359740 400 359792 406
rect 359894 354 360006 480
rect 360120 406 360148 2858
rect 360442 2802 360470 3060
rect 361546 2802 361574 3060
rect 362650 2922 362678 3060
rect 363754 2922 363782 3060
rect 362638 2916 362690 2922
rect 362638 2858 362690 2864
rect 363512 2916 363564 2922
rect 363512 2858 363564 2864
rect 363742 2916 363794 2922
rect 363742 2858 363794 2864
rect 360442 2774 360516 2802
rect 360488 678 360516 2774
rect 361500 2774 361574 2802
rect 362500 2848 362552 2854
rect 362500 2790 362552 2796
rect 360476 672 360528 678
rect 360476 614 360528 620
rect 361120 604 361172 610
rect 361120 546 361172 552
rect 361132 480 361160 546
rect 359792 348 360006 354
rect 359740 342 360006 348
rect 360108 400 360160 406
rect 360108 342 360160 348
rect 359752 326 360006 342
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361500 474 361528 2774
rect 361488 468 361540 474
rect 361488 410 361540 416
rect 362132 400 362184 406
rect 362286 354 362398 480
rect 362512 406 362540 2790
rect 363524 610 363552 2858
rect 364858 2802 364886 3060
rect 365962 2854 365990 3060
rect 366180 2916 366232 2922
rect 366180 2858 366232 2864
rect 365950 2848 366002 2854
rect 364858 2774 364932 2802
rect 365950 2790 366002 2796
rect 364904 746 364932 2774
rect 364892 740 364944 746
rect 364892 682 364944 688
rect 366192 678 366220 2858
rect 367066 2802 367094 3060
rect 367020 2774 367094 2802
rect 368170 2802 368198 3060
rect 369274 2922 369302 3060
rect 370378 2922 370406 3060
rect 369262 2916 369314 2922
rect 369262 2858 369314 2864
rect 370228 2916 370280 2922
rect 370228 2858 370280 2864
rect 370366 2916 370418 2922
rect 370366 2858 370418 2864
rect 369768 2848 369820 2854
rect 368170 2774 368336 2802
rect 369768 2790 369820 2796
rect 367020 814 367048 2774
rect 367008 808 367060 814
rect 367008 750 367060 756
rect 368308 678 368336 2774
rect 369400 740 369452 746
rect 369400 682 369452 688
rect 364616 672 364668 678
rect 364616 614 364668 620
rect 366180 672 366232 678
rect 366180 614 366232 620
rect 368204 672 368256 678
rect 368204 614 368256 620
rect 368296 672 368348 678
rect 368296 614 368348 620
rect 363512 604 363564 610
rect 363512 546 363564 552
rect 364628 480 364656 614
rect 367008 604 367060 610
rect 367008 546 367060 552
rect 367020 480 367048 546
rect 368216 480 368244 614
rect 369412 480 369440 682
rect 369780 610 369808 2790
rect 369768 604 369820 610
rect 369768 546 369820 552
rect 362184 348 362398 354
rect 362132 342 362398 348
rect 362500 400 362552 406
rect 362500 342 362552 348
rect 363482 354 363594 480
rect 363696 400 363748 406
rect 363482 348 363696 354
rect 363482 342 363748 348
rect 362144 326 362398 342
rect 362286 -960 362398 326
rect 363482 326 363736 342
rect 363482 -960 363594 326
rect 364586 -960 364698 480
rect 365628 468 365680 474
rect 365628 410 365680 416
rect 365640 354 365668 410
rect 365782 354 365894 480
rect 365640 326 365894 354
rect 365782 -960 365894 326
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370240 406 370268 2858
rect 371482 2802 371510 3060
rect 372586 2938 372614 3060
rect 372540 2910 372614 2938
rect 373690 2922 373718 3060
rect 372712 2916 372764 2922
rect 371482 2774 371556 2802
rect 370596 604 370648 610
rect 370596 546 370648 552
rect 370608 480 370636 546
rect 370228 400 370280 406
rect 370228 342 370280 348
rect 370566 -960 370678 480
rect 371528 474 371556 2774
rect 371700 808 371752 814
rect 371700 750 371752 756
rect 371712 480 371740 750
rect 371516 468 371568 474
rect 371516 410 371568 416
rect 371670 -960 371782 480
rect 372540 134 372568 2910
rect 372712 2858 372764 2864
rect 373678 2916 373730 2922
rect 373678 2858 373730 2864
rect 372724 610 372752 2858
rect 374794 2854 374822 3060
rect 375898 2922 375926 3060
rect 375104 2916 375156 2922
rect 375104 2858 375156 2864
rect 375886 2916 375938 2922
rect 375886 2858 375938 2864
rect 374782 2848 374834 2854
rect 374782 2790 374834 2796
rect 372896 672 372948 678
rect 372896 614 372948 620
rect 372712 604 372764 610
rect 372712 546 372764 552
rect 372908 480 372936 614
rect 372528 128 372580 134
rect 372528 70 372580 76
rect 372866 -960 372978 480
rect 373908 400 373960 406
rect 374062 354 374174 480
rect 375116 406 375144 2858
rect 376668 2848 376720 2854
rect 376668 2790 376720 2796
rect 377002 2802 377030 3060
rect 378106 2802 378134 3060
rect 379210 2922 379238 3060
rect 380314 2922 380342 3060
rect 378508 2916 378560 2922
rect 378508 2858 378560 2864
rect 379198 2916 379250 2922
rect 379198 2858 379250 2864
rect 380164 2916 380216 2922
rect 380164 2858 380216 2864
rect 380302 2916 380354 2922
rect 380302 2858 380354 2864
rect 376680 610 376708 2790
rect 377002 2774 377076 2802
rect 375288 604 375340 610
rect 375288 546 375340 552
rect 376668 604 376720 610
rect 376668 546 376720 552
rect 375300 480 375328 546
rect 373960 348 374174 354
rect 373908 342 374174 348
rect 375104 400 375156 406
rect 375104 342 375156 348
rect 373920 326 374174 342
rect 374062 -960 374174 326
rect 375258 -960 375370 480
rect 376300 468 376352 474
rect 376300 410 376352 416
rect 376312 354 376340 410
rect 376454 354 376566 480
rect 377048 474 377076 2774
rect 378060 2774 378134 2802
rect 378060 814 378088 2774
rect 378048 808 378100 814
rect 378048 750 378100 756
rect 378520 678 378548 2858
rect 380176 746 380204 2858
rect 381418 2802 381446 3060
rect 382280 2916 382332 2922
rect 382280 2858 382332 2864
rect 381418 2774 381492 2802
rect 380164 740 380216 746
rect 380164 682 380216 688
rect 378508 672 378560 678
rect 378508 614 378560 620
rect 381176 672 381228 678
rect 381176 614 381228 620
rect 379980 604 380032 610
rect 379980 546 380032 552
rect 379992 480 380020 546
rect 381188 480 381216 614
rect 377036 468 377088 474
rect 377036 410 377088 416
rect 376312 326 376566 354
rect 376454 -960 376566 326
rect 377650 82 377762 480
rect 378692 400 378744 406
rect 378846 354 378958 480
rect 378744 348 378958 354
rect 378692 342 378958 348
rect 378704 326 378958 342
rect 377864 128 377916 134
rect 377650 76 377864 82
rect 377650 70 377916 76
rect 377650 54 377904 70
rect 377650 -960 377762 54
rect 378846 -960 378958 326
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 381464 202 381492 2774
rect 382292 610 382320 2858
rect 382522 2854 382550 3060
rect 382510 2848 382562 2854
rect 383626 2802 383654 3060
rect 384730 2802 384758 3060
rect 382510 2790 382562 2796
rect 383396 2774 383654 2802
rect 384684 2774 384758 2802
rect 385834 2802 385862 3060
rect 386938 2922 386966 3060
rect 388042 2922 388070 3060
rect 386926 2916 386978 2922
rect 386926 2858 386978 2864
rect 387892 2916 387944 2922
rect 387892 2858 387944 2864
rect 388030 2916 388082 2922
rect 388030 2858 388082 2864
rect 387708 2848 387760 2854
rect 385834 2774 385908 2802
rect 387708 2790 387760 2796
rect 382280 604 382332 610
rect 382280 546 382332 552
rect 382188 468 382240 474
rect 382188 410 382240 416
rect 382200 354 382228 410
rect 382342 354 382454 480
rect 382200 326 382454 354
rect 381452 196 381504 202
rect 381452 138 381504 144
rect 382342 -960 382454 326
rect 383396 134 383424 2774
rect 383568 808 383620 814
rect 383568 750 383620 756
rect 383580 480 383608 750
rect 384684 678 384712 2774
rect 385880 814 385908 2774
rect 385868 808 385920 814
rect 385868 750 385920 756
rect 384764 740 384816 746
rect 384764 682 384816 688
rect 384672 672 384724 678
rect 384672 614 384724 620
rect 384776 480 384804 682
rect 385960 604 386012 610
rect 385960 546 386012 552
rect 385972 480 386000 546
rect 383384 128 383436 134
rect 383384 70 383436 76
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 218 387238 480
rect 387720 354 387748 2790
rect 387904 474 387932 2858
rect 389146 2802 389174 3060
rect 389100 2774 389174 2802
rect 390250 2802 390278 3060
rect 391354 2922 391382 3060
rect 390652 2916 390704 2922
rect 390652 2858 390704 2864
rect 391342 2916 391394 2922
rect 391342 2858 391394 2864
rect 390250 2774 390324 2802
rect 389100 678 389128 2774
rect 389088 672 389140 678
rect 389088 614 389140 620
rect 387892 468 387944 474
rect 387892 410 387944 416
rect 388230 354 388342 480
rect 387720 326 388342 354
rect 386984 202 387238 218
rect 386972 196 387238 202
rect 387024 190 387238 196
rect 386972 138 387024 144
rect 387126 -960 387238 190
rect 388230 -960 388342 326
rect 389426 82 389538 480
rect 390296 270 390324 2774
rect 390664 746 390692 2858
rect 392458 2802 392486 3060
rect 393562 2854 393590 3060
rect 394666 2938 394694 3060
rect 394424 2916 394476 2922
rect 394424 2858 394476 2864
rect 394528 2910 394694 2938
rect 393550 2848 393602 2854
rect 392458 2774 392532 2802
rect 393550 2790 393602 2796
rect 391848 808 391900 814
rect 391848 750 391900 756
rect 390652 740 390704 746
rect 390652 682 390704 688
rect 390652 604 390704 610
rect 390652 546 390704 552
rect 390664 480 390692 546
rect 391860 480 391888 750
rect 390284 264 390336 270
rect 390284 206 390336 212
rect 389640 128 389692 134
rect 389426 76 389640 82
rect 389426 70 389692 76
rect 389426 54 389680 70
rect 389426 -960 389538 54
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392504 406 392532 2774
rect 394240 740 394292 746
rect 394240 682 394292 688
rect 394252 480 394280 682
rect 394436 610 394464 2858
rect 394528 814 394556 2910
rect 395770 2802 395798 3060
rect 396874 2922 396902 3060
rect 396862 2916 396914 2922
rect 396862 2858 396914 2864
rect 397978 2854 398006 3060
rect 399082 2922 399110 3060
rect 398748 2916 398800 2922
rect 398748 2858 398800 2864
rect 399070 2916 399122 2922
rect 399070 2858 399122 2864
rect 396724 2848 396776 2854
rect 395770 2774 395844 2802
rect 396724 2790 396776 2796
rect 397966 2848 398018 2854
rect 397966 2790 398018 2796
rect 394516 808 394568 814
rect 394516 750 394568 756
rect 395816 678 395844 2774
rect 396736 746 396764 2790
rect 396724 740 396776 746
rect 396724 682 396776 688
rect 398760 678 398788 2858
rect 399852 2848 399904 2854
rect 400186 2802 400214 3060
rect 399852 2790 399904 2796
rect 395344 672 395396 678
rect 395344 614 395396 620
rect 395804 672 395856 678
rect 395804 614 395856 620
rect 398748 672 398800 678
rect 398748 614 398800 620
rect 394424 604 394476 610
rect 394424 546 394476 552
rect 395356 480 395384 614
rect 397736 604 397788 610
rect 397736 546 397788 552
rect 397748 480 397776 546
rect 392860 468 392912 474
rect 392860 410 392912 416
rect 392492 400 392544 406
rect 392492 342 392544 348
rect 392872 354 392900 410
rect 393014 354 393126 480
rect 392872 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396356 264 396408 270
rect 396510 218 396622 480
rect 396408 212 396622 218
rect 396356 206 396622 212
rect 396368 190 396622 206
rect 396510 -960 396622 190
rect 397706 -960 397818 480
rect 398748 400 398800 406
rect 398902 354 399014 480
rect 399864 406 399892 2790
rect 399956 2774 400214 2802
rect 401290 2802 401318 3060
rect 402394 2922 402422 3060
rect 401600 2916 401652 2922
rect 401600 2858 401652 2864
rect 402382 2916 402434 2922
rect 402382 2858 402434 2864
rect 401290 2774 401548 2802
rect 398800 348 399014 354
rect 398748 342 399014 348
rect 399852 400 399904 406
rect 399852 342 399904 348
rect 398760 326 399014 342
rect 398902 -960 399014 326
rect 399956 202 399984 2774
rect 401324 808 401376 814
rect 401324 750 401376 756
rect 400128 740 400180 746
rect 400128 682 400180 688
rect 400140 480 400168 682
rect 401336 480 401364 750
rect 399944 196 399996 202
rect 399944 138 399996 144
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 401520 270 401548 2774
rect 401612 542 401640 2858
rect 403498 2854 403526 3060
rect 404268 2916 404320 2922
rect 404268 2858 404320 2864
rect 403486 2848 403538 2854
rect 403486 2790 403538 2796
rect 403624 672 403676 678
rect 403624 614 403676 620
rect 402520 604 402572 610
rect 402520 546 402572 552
rect 401600 536 401652 542
rect 401600 478 401652 484
rect 402532 480 402560 546
rect 403636 480 403664 614
rect 401508 264 401560 270
rect 401508 206 401560 212
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404280 338 404308 2858
rect 404602 2802 404630 3060
rect 405706 2802 405734 3060
rect 406810 2922 406838 3060
rect 407914 2922 407942 3060
rect 406798 2916 406850 2922
rect 406798 2858 406850 2864
rect 407764 2916 407816 2922
rect 407764 2858 407816 2864
rect 407902 2916 407954 2922
rect 407902 2858 407954 2864
rect 404602 2774 404676 2802
rect 404648 814 404676 2774
rect 405660 2774 405734 2802
rect 407028 2848 407080 2854
rect 407028 2790 407080 2796
rect 404636 808 404688 814
rect 404636 750 404688 756
rect 404636 400 404688 406
rect 404790 354 404902 480
rect 404688 348 404902 354
rect 404636 342 404902 348
rect 404268 332 404320 338
rect 404648 326 404902 342
rect 404268 274 404320 280
rect 404790 -960 404902 326
rect 405660 134 405688 2774
rect 407040 678 407068 2790
rect 407776 746 407804 2858
rect 409018 2854 409046 3060
rect 409788 2916 409840 2922
rect 409788 2858 409840 2864
rect 409006 2848 409058 2854
rect 409006 2790 409058 2796
rect 407764 740 407816 746
rect 407764 682 407816 688
rect 407028 672 407080 678
rect 407028 614 407080 620
rect 409800 610 409828 2858
rect 410122 2802 410150 3060
rect 411226 2802 411254 3060
rect 410122 2774 410196 2802
rect 406016 604 406068 610
rect 406016 546 406068 552
rect 409788 604 409840 610
rect 409788 546 409840 552
rect 406028 480 406056 546
rect 405648 128 405700 134
rect 405648 70 405700 76
rect 405986 -960 406098 480
rect 407182 218 407294 480
rect 407040 202 407294 218
rect 407028 196 407294 202
rect 407080 190 407294 196
rect 407028 138 407080 144
rect 407182 -960 407294 190
rect 408378 218 408490 480
rect 409574 354 409686 480
rect 409432 338 409686 354
rect 410168 338 410196 2774
rect 411180 2774 411254 2802
rect 412330 2802 412358 3060
rect 413434 2802 413462 3060
rect 414538 2802 414566 3060
rect 415642 2922 415670 3060
rect 415630 2916 415682 2922
rect 415630 2858 415682 2864
rect 416596 2848 416648 2854
rect 412330 2774 412404 2802
rect 413434 2774 413508 2802
rect 414538 2774 414612 2802
rect 416746 2802 416774 3060
rect 417850 2802 417878 3060
rect 416596 2790 416648 2796
rect 410800 672 410852 678
rect 410800 614 410852 620
rect 410812 480 410840 614
rect 409420 332 409686 338
rect 409472 326 409686 332
rect 409420 274 409472 280
rect 408592 264 408644 270
rect 408378 212 408592 218
rect 408378 206 408644 212
rect 408378 190 408632 206
rect 408378 -960 408490 190
rect 409574 -960 409686 326
rect 410156 332 410208 338
rect 410156 274 410208 280
rect 410770 -960 410882 480
rect 411180 202 411208 2774
rect 411904 808 411956 814
rect 411904 750 411956 756
rect 411916 480 411944 750
rect 411168 196 411220 202
rect 411168 138 411220 144
rect 411874 -960 411986 480
rect 412376 270 412404 2774
rect 412364 264 412416 270
rect 412364 206 412416 212
rect 412916 128 412968 134
rect 413070 82 413182 480
rect 413480 134 413508 2774
rect 414584 746 414612 2774
rect 414296 740 414348 746
rect 414296 682 414348 688
rect 414572 740 414624 746
rect 414572 682 414624 688
rect 414308 480 414336 682
rect 416608 626 416636 2790
rect 416700 2774 416774 2802
rect 417804 2774 417878 2802
rect 418954 2802 418982 3060
rect 420058 2802 420086 3060
rect 418954 2774 419212 2802
rect 416700 814 416728 2774
rect 416688 808 416740 814
rect 416688 750 416740 756
rect 417804 678 417832 2774
rect 417792 672 417844 678
rect 415492 604 415544 610
rect 416608 598 416728 626
rect 417792 614 417844 620
rect 415492 546 415544 552
rect 415504 480 415532 546
rect 416700 480 416728 598
rect 417884 604 417936 610
rect 417884 546 417936 552
rect 418816 598 419028 626
rect 417896 480 417924 546
rect 412968 76 413182 82
rect 412916 70 413182 76
rect 413468 128 413520 134
rect 413468 70 413520 76
rect 412928 54 413182 70
rect 413070 -960 413182 54
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418816 202 418844 598
rect 419000 480 419028 598
rect 418804 196 418856 202
rect 418804 138 418856 144
rect 418958 -960 419070 480
rect 419184 406 419212 2774
rect 420012 2774 420086 2802
rect 421162 2802 421190 3060
rect 422266 2904 422294 3060
rect 422266 2876 422340 2904
rect 422312 2802 422340 2876
rect 421162 2774 421236 2802
rect 420012 474 420040 2774
rect 421208 610 421236 2774
rect 422220 2774 422340 2802
rect 423370 2802 423398 3060
rect 424474 2922 424502 3060
rect 425578 2922 425606 3060
rect 423772 2916 423824 2922
rect 423772 2858 423824 2864
rect 424462 2916 424514 2922
rect 424462 2858 424514 2864
rect 425428 2916 425480 2922
rect 425428 2858 425480 2864
rect 425566 2916 425618 2922
rect 425566 2858 425618 2864
rect 423370 2774 423444 2802
rect 421196 604 421248 610
rect 421196 546 421248 552
rect 420000 468 420052 474
rect 420000 410 420052 416
rect 419172 400 419224 406
rect 419172 342 419224 348
rect 420154 218 420266 480
rect 420368 264 420420 270
rect 420154 212 420368 218
rect 420154 206 420420 212
rect 420154 190 420408 206
rect 420154 -960 420266 190
rect 421196 128 421248 134
rect 421350 82 421462 480
rect 422220 202 422248 2774
rect 422576 740 422628 746
rect 422576 682 422628 688
rect 422588 480 422616 682
rect 422208 196 422260 202
rect 422208 138 422260 144
rect 421248 76 421462 82
rect 421196 70 421462 76
rect 421208 54 421462 70
rect 421350 -960 421462 54
rect 422546 -960 422658 480
rect 423416 270 423444 2774
rect 423784 480 423812 2858
rect 424968 808 425020 814
rect 424968 750 425020 756
rect 424980 480 425008 750
rect 425440 746 425468 2858
rect 426682 2802 426710 3060
rect 427786 2802 427814 3060
rect 428890 2922 428918 3060
rect 429994 2922 430022 3060
rect 428740 2916 428792 2922
rect 428740 2858 428792 2864
rect 428878 2916 428930 2922
rect 428878 2858 428930 2864
rect 429844 2916 429896 2922
rect 429844 2858 429896 2864
rect 429982 2916 430034 2922
rect 429982 2858 430034 2864
rect 426682 2774 426756 2802
rect 425428 740 425480 746
rect 425428 682 425480 688
rect 423404 264 423456 270
rect 423404 206 423456 212
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 354 426246 480
rect 425992 338 426246 354
rect 426728 338 426756 2774
rect 427740 2774 427814 2802
rect 427084 400 427136 406
rect 427238 354 427350 480
rect 427136 348 427350 354
rect 427084 342 427350 348
rect 425980 332 426246 338
rect 426032 326 426246 332
rect 425980 274 426032 280
rect 426134 -960 426246 326
rect 426716 332 426768 338
rect 427096 326 427350 342
rect 426716 274 426768 280
rect 427238 -960 427350 326
rect 427740 134 427768 2774
rect 428752 678 428780 2858
rect 428740 672 428792 678
rect 428740 614 428792 620
rect 429660 604 429712 610
rect 429660 546 429712 552
rect 429672 480 429700 546
rect 428434 354 428546 480
rect 428648 468 428700 474
rect 428648 410 428700 416
rect 428660 354 428688 410
rect 428434 326 428688 354
rect 427728 128 427780 134
rect 427728 70 427780 76
rect 428434 -960 428546 326
rect 429630 -960 429742 480
rect 429856 474 429884 2858
rect 431098 2802 431126 3060
rect 432202 2854 432230 3060
rect 433156 2916 433208 2922
rect 433156 2858 433208 2864
rect 432190 2848 432242 2854
rect 431098 2774 431172 2802
rect 432190 2790 432242 2796
rect 429844 468 429896 474
rect 429844 410 429896 416
rect 430826 218 430938 480
rect 431144 338 431172 2774
rect 433064 876 433116 882
rect 433064 818 433116 824
rect 431132 332 431184 338
rect 431132 274 431184 280
rect 431868 264 431920 270
rect 430826 202 431080 218
rect 432022 218 432134 480
rect 431920 212 432134 218
rect 431868 206 432134 212
rect 430826 196 431092 202
rect 430826 190 431040 196
rect 430826 -960 430938 190
rect 431880 190 432134 206
rect 433076 202 433104 818
rect 433168 814 433196 2858
rect 433306 2802 433334 3060
rect 433260 2774 433334 2802
rect 434410 2802 434438 3060
rect 435514 2802 435542 3060
rect 436618 2802 436646 3060
rect 434410 2774 434668 2802
rect 435514 2774 435772 2802
rect 433260 882 433288 2774
rect 433248 876 433300 882
rect 433248 818 433300 824
rect 433156 808 433208 814
rect 433156 750 433208 756
rect 433248 740 433300 746
rect 433248 682 433300 688
rect 433260 480 433288 682
rect 434444 672 434496 678
rect 434444 614 434496 620
rect 434456 480 434484 614
rect 431040 138 431092 144
rect 432022 -960 432134 190
rect 433064 196 433116 202
rect 433064 138 433116 144
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 434640 270 434668 2774
rect 435548 604 435600 610
rect 435548 546 435600 552
rect 435560 480 435588 546
rect 434628 264 434680 270
rect 434628 206 434680 212
rect 435518 -960 435630 480
rect 435744 406 435772 2774
rect 436572 2774 436646 2802
rect 437722 2802 437750 3060
rect 438826 2802 438854 3060
rect 439930 2922 439958 3060
rect 439918 2916 439970 2922
rect 439918 2858 439970 2864
rect 437722 2774 437796 2802
rect 436572 542 436600 2774
rect 437768 610 437796 2774
rect 438780 2774 438854 2802
rect 438952 2848 439004 2854
rect 438952 2790 439004 2796
rect 441034 2802 441062 3060
rect 442138 2854 442166 3060
rect 442908 2916 442960 2922
rect 442908 2858 442960 2864
rect 442126 2848 442178 2854
rect 437940 672 437992 678
rect 437940 614 437992 620
rect 437756 604 437808 610
rect 437756 546 437808 552
rect 436560 536 436612 542
rect 436560 478 436612 484
rect 437952 480 437980 614
rect 435732 400 435784 406
rect 435732 342 435784 348
rect 436714 82 436826 480
rect 436928 128 436980 134
rect 436714 76 436928 82
rect 436714 70 436980 76
rect 436714 54 436968 70
rect 436714 -960 436826 54
rect 437910 -960 438022 480
rect 438780 134 438808 2774
rect 438964 678 438992 2790
rect 441034 2774 441108 2802
rect 442126 2790 442178 2796
rect 439136 808 439188 814
rect 439136 750 439188 756
rect 438952 672 439004 678
rect 438952 614 439004 620
rect 439148 480 439176 750
rect 438768 128 438820 134
rect 438768 70 438820 76
rect 439106 -960 439218 480
rect 440302 354 440414 480
rect 440160 338 440414 354
rect 441080 338 441108 2774
rect 442920 678 442948 2858
rect 443242 2802 443270 3060
rect 444346 2802 444374 3060
rect 443242 2774 443316 2802
rect 443288 814 443316 2774
rect 444300 2774 444374 2802
rect 445450 2802 445478 3060
rect 446554 2802 446582 3060
rect 447658 2802 447686 3060
rect 448762 2802 448790 3060
rect 449866 2802 449894 3060
rect 450970 2922 450998 3060
rect 450958 2916 451010 2922
rect 450958 2858 451010 2864
rect 452074 2854 452102 3060
rect 452568 2916 452620 2922
rect 452568 2858 452620 2864
rect 445450 2774 445524 2802
rect 446554 2774 446628 2802
rect 447658 2774 447732 2802
rect 448762 2774 448836 2802
rect 443276 808 443328 814
rect 443276 750 443328 756
rect 441528 672 441580 678
rect 441528 614 441580 620
rect 442908 672 442960 678
rect 442908 614 442960 620
rect 441540 480 441568 614
rect 440148 332 440414 338
rect 440200 326 440414 332
rect 440148 274 440200 280
rect 440302 -960 440414 326
rect 441068 332 441120 338
rect 441068 274 441120 280
rect 441498 -960 441610 480
rect 442602 218 442714 480
rect 443644 264 443696 270
rect 442602 202 442856 218
rect 443798 218 443910 480
rect 443696 212 443910 218
rect 443644 206 443910 212
rect 442602 196 442868 202
rect 442602 190 442816 196
rect 442602 -960 442714 190
rect 443656 190 443910 206
rect 444300 202 444328 2774
rect 444994 354 445106 480
rect 445208 400 445260 406
rect 444994 348 445208 354
rect 444994 342 445260 348
rect 444994 326 445248 342
rect 442816 138 442868 144
rect 443798 -960 443910 190
rect 444288 196 444340 202
rect 444288 138 444340 144
rect 444994 -960 445106 326
rect 445496 270 445524 2774
rect 446036 536 446088 542
rect 446036 478 446088 484
rect 446048 354 446076 478
rect 446190 354 446302 480
rect 446600 406 446628 2774
rect 447704 678 447732 2774
rect 448808 746 448836 2774
rect 449636 2774 449894 2802
rect 451188 2848 451240 2854
rect 451188 2790 451240 2796
rect 452062 2848 452114 2854
rect 452062 2790 452114 2796
rect 448796 740 448848 746
rect 448796 682 448848 688
rect 447692 672 447744 678
rect 447692 614 447744 620
rect 447416 604 447468 610
rect 447416 546 447468 552
rect 447428 480 447456 546
rect 446048 326 446302 354
rect 446588 400 446640 406
rect 446588 342 446640 348
rect 445484 264 445536 270
rect 445484 206 445536 212
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448428 128 448480 134
rect 448582 82 448694 480
rect 449636 134 449664 2774
rect 451096 808 451148 814
rect 451096 750 451148 756
rect 449808 604 449860 610
rect 449808 546 449860 552
rect 450912 604 450964 610
rect 450912 546 450964 552
rect 449820 480 449848 546
rect 450924 480 450952 546
rect 448480 76 448694 82
rect 448428 70 448694 76
rect 449624 128 449676 134
rect 449624 70 449676 76
rect 448440 54 448694 70
rect 448582 -960 448694 54
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451108 474 451136 750
rect 451200 610 451228 2790
rect 452580 610 452608 2858
rect 453178 2802 453206 3060
rect 453132 2774 453206 2802
rect 454282 2802 454310 3060
rect 455386 2802 455414 3060
rect 454282 2774 454356 2802
rect 451188 604 451240 610
rect 451188 546 451240 552
rect 452108 604 452160 610
rect 452108 546 452160 552
rect 452568 604 452620 610
rect 452568 546 452620 552
rect 452120 480 452148 546
rect 451096 468 451148 474
rect 451096 410 451148 416
rect 452078 -960 452190 480
rect 453132 338 453160 2774
rect 454328 542 454356 2774
rect 455340 2774 455414 2802
rect 456490 2802 456518 3060
rect 457594 2802 457622 3060
rect 458698 2802 458726 3060
rect 459802 2802 459830 3060
rect 460906 2802 460934 3060
rect 462010 2922 462038 3060
rect 463114 2922 463142 3060
rect 464218 2922 464246 3060
rect 461998 2916 462050 2922
rect 461998 2858 462050 2864
rect 463102 2916 463154 2922
rect 463102 2858 463154 2864
rect 464068 2916 464120 2922
rect 464068 2858 464120 2864
rect 464206 2916 464258 2922
rect 464206 2858 464258 2864
rect 456490 2774 456564 2802
rect 457594 2774 457668 2802
rect 458698 2774 458772 2802
rect 459802 2774 459876 2802
rect 454316 536 454368 542
rect 453274 354 453386 480
rect 454316 478 454368 484
rect 453488 468 453540 474
rect 453488 410 453540 416
rect 453500 354 453528 410
rect 453120 332 453172 338
rect 453120 274 453172 280
rect 453274 326 453528 354
rect 453274 -960 453386 326
rect 454470 218 454582 480
rect 454328 202 454582 218
rect 455340 202 455368 2774
rect 455666 218 455778 480
rect 456536 270 456564 2774
rect 456708 400 456760 406
rect 456862 354 456974 480
rect 457640 474 457668 2774
rect 458744 678 458772 2774
rect 459848 746 459876 2774
rect 460860 2774 460934 2802
rect 462228 2848 462280 2854
rect 462228 2790 462280 2796
rect 463608 2848 463660 2854
rect 463608 2790 463660 2796
rect 459192 740 459244 746
rect 459192 682 459244 688
rect 459836 740 459888 746
rect 459836 682 459888 688
rect 458088 672 458140 678
rect 458088 614 458140 620
rect 458732 672 458784 678
rect 458732 614 458784 620
rect 458100 480 458128 614
rect 459204 480 459232 682
rect 457628 468 457680 474
rect 457628 410 457680 416
rect 456760 348 456974 354
rect 456708 342 456974 348
rect 456720 326 456974 342
rect 455880 264 455932 270
rect 455666 212 455880 218
rect 455666 206 455932 212
rect 456524 264 456576 270
rect 456524 206 456576 212
rect 454316 196 454582 202
rect 454368 190 454582 196
rect 454316 138 454368 144
rect 454470 -960 454582 190
rect 455328 196 455380 202
rect 455328 138 455380 144
rect 455666 190 455920 206
rect 455666 -960 455778 190
rect 456862 -960 456974 326
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460204 128 460256 134
rect 460358 82 460470 480
rect 460860 134 460888 2774
rect 461584 604 461636 610
rect 461584 546 461636 552
rect 461596 480 461624 546
rect 460256 76 460470 82
rect 460204 70 460470 76
rect 460848 128 460900 134
rect 460848 70 460900 76
rect 460216 54 460470 70
rect 460358 -960 460470 54
rect 461554 -960 461666 480
rect 462240 354 462268 2790
rect 463620 746 463648 2790
rect 464080 882 464108 2858
rect 465322 2854 465350 3060
rect 466426 2938 466454 3060
rect 466184 2916 466236 2922
rect 466184 2858 466236 2864
rect 466288 2910 466454 2938
rect 465310 2848 465362 2854
rect 465310 2790 465362 2796
rect 466196 950 466224 2858
rect 466184 944 466236 950
rect 466184 886 466236 892
rect 464068 876 464120 882
rect 464068 818 464120 824
rect 463608 740 463660 746
rect 463608 682 463660 688
rect 466288 626 466316 2910
rect 467530 2802 467558 3060
rect 468634 2802 468662 3060
rect 469738 2802 469766 3060
rect 470842 2802 470870 3060
rect 471946 2802 471974 3060
rect 467530 2774 467696 2802
rect 468634 2774 468892 2802
rect 469738 2774 469812 2802
rect 470842 2774 470916 2802
rect 467288 672 467340 678
rect 466288 598 466500 626
rect 467288 614 467340 620
rect 464988 536 465040 542
rect 462750 354 462862 480
rect 462240 326 462862 354
rect 462750 -960 462862 326
rect 463946 354 464058 480
rect 464988 478 465040 484
rect 465000 354 465028 478
rect 465142 354 465254 480
rect 463946 338 464200 354
rect 463946 332 464212 338
rect 463946 326 464160 332
rect 463946 -960 464058 326
rect 465000 326 465254 354
rect 464160 274 464212 280
rect 465142 -960 465254 326
rect 466246 218 466358 480
rect 466104 202 466358 218
rect 466472 202 466500 598
rect 466092 196 466358 202
rect 466144 190 466358 196
rect 466092 138 466144 144
rect 466246 -960 466358 190
rect 466460 196 466512 202
rect 466460 138 466512 144
rect 467300 66 467328 614
rect 467472 604 467524 610
rect 467472 546 467524 552
rect 467484 480 467512 546
rect 467288 60 467340 66
rect 467288 2 467340 8
rect 467442 -960 467554 480
rect 467668 406 467696 2774
rect 468576 672 468628 678
rect 468628 620 468708 626
rect 468576 614 468708 620
rect 468588 598 468708 614
rect 468680 480 468708 598
rect 468864 542 468892 2774
rect 469784 678 469812 2774
rect 470888 1018 470916 2774
rect 471900 2774 471974 2802
rect 473050 2802 473078 3060
rect 474154 2802 474182 3060
rect 475258 2802 475286 3060
rect 476362 2922 476390 3060
rect 476350 2916 476402 2922
rect 476350 2858 476402 2864
rect 476948 2848 477000 2854
rect 473050 2774 473124 2802
rect 474154 2774 474228 2802
rect 475258 2774 475332 2802
rect 477466 2802 477494 3060
rect 478328 2916 478380 2922
rect 478328 2858 478380 2864
rect 476948 2790 477000 2796
rect 470876 1012 470928 1018
rect 470876 954 470928 960
rect 471060 808 471112 814
rect 471060 750 471112 756
rect 469772 672 469824 678
rect 469772 614 469824 620
rect 468852 536 468904 542
rect 467656 400 467708 406
rect 467656 342 467708 348
rect 468638 -960 468750 480
rect 468852 478 468904 484
rect 471072 480 471100 750
rect 469834 82 469946 480
rect 469834 66 470088 82
rect 469834 60 470100 66
rect 469834 54 470048 60
rect 469834 -960 469946 54
rect 470048 2 470100 8
rect 471030 -960 471142 480
rect 471900 270 471928 2774
rect 471888 264 471940 270
rect 471888 206 471940 212
rect 472226 82 472338 480
rect 473096 338 473124 2774
rect 474200 610 474228 2774
rect 475304 882 475332 2774
rect 475752 944 475804 950
rect 475752 886 475804 892
rect 474556 876 474608 882
rect 474556 818 474608 824
rect 475292 876 475344 882
rect 475292 818 475344 824
rect 473452 604 473504 610
rect 473452 546 473504 552
rect 474188 604 474240 610
rect 474188 546 474240 552
rect 473464 480 473492 546
rect 474568 480 474596 818
rect 475764 480 475792 886
rect 476960 480 476988 2790
rect 477420 2774 477494 2802
rect 473084 332 473136 338
rect 473084 274 473136 280
rect 472440 128 472492 134
rect 472226 76 472440 82
rect 472226 70 472492 76
rect 472226 54 472480 70
rect 472226 -960 472338 54
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 477420 134 477448 2774
rect 478340 950 478368 2858
rect 478570 2854 478598 3060
rect 478558 2848 478610 2854
rect 478558 2790 478610 2796
rect 479674 2802 479702 3060
rect 480778 2802 480806 3060
rect 481882 2802 481910 3060
rect 482986 2802 483014 3060
rect 479674 2774 479748 2802
rect 480778 2774 480852 2802
rect 481882 2774 481956 2802
rect 478328 944 478380 950
rect 478328 886 478380 892
rect 478114 218 478226 480
rect 479156 400 479208 406
rect 479310 354 479422 480
rect 479720 474 479748 2774
rect 480824 746 480852 2774
rect 481928 814 481956 2774
rect 482940 2774 483014 2802
rect 484090 2802 484118 3060
rect 485194 2802 485222 3060
rect 486298 2802 486326 3060
rect 487402 2802 487430 3060
rect 488506 2802 488534 3060
rect 484090 2774 484256 2802
rect 485194 2774 485360 2802
rect 486298 2774 486372 2802
rect 487402 2774 487476 2802
rect 482836 1012 482888 1018
rect 482836 954 482888 960
rect 481916 808 481968 814
rect 481916 750 481968 756
rect 480812 740 480864 746
rect 480812 682 480864 688
rect 481732 672 481784 678
rect 481732 614 481784 620
rect 480720 536 480772 542
rect 479708 468 479760 474
rect 479708 410 479760 416
rect 479208 348 479422 354
rect 479156 342 479422 348
rect 479168 326 479422 342
rect 478114 202 478368 218
rect 478114 196 478380 202
rect 478114 190 478328 196
rect 477408 128 477460 134
rect 477408 70 477460 76
rect 478114 -960 478226 190
rect 478328 138 478380 144
rect 479310 -960 479422 326
rect 480506 354 480618 480
rect 480720 478 480772 484
rect 481744 480 481772 614
rect 482848 480 482876 954
rect 482940 678 482968 2774
rect 482928 672 482980 678
rect 482928 614 482980 620
rect 483860 598 484072 626
rect 480732 354 480760 478
rect 480506 326 480760 354
rect 480506 -960 480618 326
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 483860 270 483888 598
rect 484044 480 484072 598
rect 483848 264 483900 270
rect 483848 206 483900 212
rect 484002 -960 484114 480
rect 484228 406 484256 2774
rect 485332 2746 485452 2774
rect 485056 598 485268 626
rect 484216 400 484268 406
rect 484216 342 484268 348
rect 485056 338 485084 598
rect 485240 480 485268 598
rect 485424 542 485452 2746
rect 486344 678 486372 2774
rect 487448 1018 487476 2774
rect 488460 2774 488534 2802
rect 488632 2848 488684 2854
rect 488632 2790 488684 2796
rect 489610 2802 489638 3060
rect 490714 2922 490742 3060
rect 490702 2916 490754 2922
rect 490702 2858 490754 2864
rect 491818 2854 491846 3060
rect 492588 2916 492640 2922
rect 492588 2858 492640 2864
rect 491806 2848 491858 2854
rect 487436 1012 487488 1018
rect 487436 954 487488 960
rect 487620 876 487672 882
rect 487620 818 487672 824
rect 485504 672 485556 678
rect 485504 614 485556 620
rect 486332 672 486384 678
rect 486332 614 486384 620
rect 485412 536 485464 542
rect 485044 332 485096 338
rect 485044 274 485096 280
rect 485198 -960 485310 480
rect 485412 478 485464 484
rect 485516 338 485544 614
rect 486424 604 486476 610
rect 486424 546 486476 552
rect 486436 480 486464 546
rect 487632 480 487660 818
rect 485504 332 485556 338
rect 485504 274 485556 280
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488460 270 488488 2774
rect 488448 264 488500 270
rect 488448 206 488500 212
rect 488644 202 488672 2790
rect 489610 2774 489684 2802
rect 491806 2790 491858 2796
rect 488816 944 488868 950
rect 488816 886 488868 892
rect 488828 480 488856 886
rect 489656 610 489684 2774
rect 492600 950 492628 2858
rect 492922 2802 492950 3060
rect 494026 2802 494054 3060
rect 492922 2774 492996 2802
rect 492588 944 492640 950
rect 492588 886 492640 892
rect 492968 882 492996 2774
rect 493980 2774 494054 2802
rect 495130 2802 495158 3060
rect 496234 2802 496262 3060
rect 497338 2802 497366 3060
rect 498442 2802 498470 3060
rect 499546 2802 499574 3060
rect 495130 2774 495204 2802
rect 496234 2774 496308 2802
rect 497338 2774 497412 2802
rect 498442 2774 498516 2802
rect 492956 876 493008 882
rect 492956 818 493008 824
rect 493508 740 493560 746
rect 493508 682 493560 688
rect 489644 604 489696 610
rect 489644 546 489696 552
rect 493520 480 493548 682
rect 488632 196 488684 202
rect 488632 138 488684 144
rect 488786 -960 488898 480
rect 489890 82 490002 480
rect 491086 218 491198 480
rect 490944 202 491198 218
rect 490932 196 491198 202
rect 490984 190 491198 196
rect 490932 138 490984 144
rect 490104 128 490156 134
rect 489890 76 490104 82
rect 489890 70 490156 76
rect 489890 54 490144 70
rect 489890 -960 490002 54
rect 491086 -960 491198 190
rect 492282 354 492394 480
rect 492496 468 492548 474
rect 492496 410 492548 416
rect 492508 354 492536 410
rect 492282 326 492536 354
rect 492282 -960 492394 326
rect 493478 -960 493590 480
rect 493980 134 494008 2774
rect 494704 808 494756 814
rect 494704 750 494756 756
rect 494716 480 494744 750
rect 493968 128 494020 134
rect 493968 70 494020 76
rect 494674 -960 494786 480
rect 495176 202 495204 2774
rect 495870 354 495982 480
rect 496280 474 496308 2774
rect 497384 678 497412 2774
rect 498488 814 498516 2774
rect 499500 2774 499574 2802
rect 500650 2802 500678 3060
rect 501754 2802 501782 3060
rect 502858 2802 502886 3060
rect 500650 2774 500816 2802
rect 501754 2774 501828 2802
rect 498476 808 498528 814
rect 498476 750 498528 756
rect 499396 740 499448 746
rect 499396 682 499448 688
rect 497372 672 497424 678
rect 497372 614 497424 620
rect 498384 536 498436 542
rect 496268 468 496320 474
rect 496268 410 496320 416
rect 495728 338 495982 354
rect 495716 332 495982 338
rect 495768 326 495982 332
rect 495716 274 495768 280
rect 495164 196 495216 202
rect 495164 138 495216 144
rect 495870 -960 495982 326
rect 497066 354 497178 480
rect 497280 400 497332 406
rect 497066 348 497280 354
rect 497066 342 497332 348
rect 498170 354 498282 480
rect 498384 478 498436 484
rect 499408 480 499436 682
rect 499500 626 499528 2774
rect 500592 1012 500644 1018
rect 500592 954 500644 960
rect 499500 598 499620 626
rect 498396 354 498424 478
rect 497066 326 497320 342
rect 498170 326 498424 354
rect 497066 -960 497178 326
rect 498170 -960 498282 326
rect 499366 -960 499478 480
rect 499592 338 499620 598
rect 500604 480 500632 954
rect 499580 332 499632 338
rect 499580 274 499632 280
rect 500562 -960 500674 480
rect 500788 406 500816 2774
rect 501800 1018 501828 2774
rect 502812 2774 502886 2802
rect 503962 2802 503990 3060
rect 505066 2802 505094 3060
rect 506170 2922 506198 3060
rect 506158 2916 506210 2922
rect 506158 2858 506210 2864
rect 503962 2774 504036 2802
rect 501788 1012 501840 1018
rect 501788 954 501840 960
rect 501616 598 501828 626
rect 500776 400 500828 406
rect 500776 342 500828 348
rect 501616 270 501644 598
rect 501800 480 501828 598
rect 502812 542 502840 2774
rect 504008 950 504036 2774
rect 505020 2774 505094 2802
rect 505376 2848 505428 2854
rect 505376 2790 505428 2796
rect 507274 2802 507302 3060
rect 508378 2922 508406 3060
rect 507860 2916 507912 2922
rect 507860 2858 507912 2864
rect 508366 2916 508418 2922
rect 508366 2858 508418 2864
rect 503996 944 504048 950
rect 503996 886 504048 892
rect 504180 876 504232 882
rect 504180 818 504232 824
rect 503628 808 503680 814
rect 503904 808 503956 814
rect 503680 756 503904 762
rect 503628 750 503956 756
rect 503640 734 503944 750
rect 502984 604 503036 610
rect 502984 546 503036 552
rect 502800 536 502852 542
rect 501604 264 501656 270
rect 501604 206 501656 212
rect 501758 -960 501870 480
rect 502800 478 502852 484
rect 502996 480 503024 546
rect 504192 480 504220 818
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505020 270 505048 2774
rect 505388 480 505416 2790
rect 507274 2774 507348 2802
rect 506112 1012 506164 1018
rect 506112 954 506164 960
rect 506124 542 506152 954
rect 507320 882 507348 2774
rect 507872 1018 507900 2858
rect 509482 2854 509510 3060
rect 509976 2916 510028 2922
rect 509976 2858 510028 2864
rect 509470 2848 509522 2854
rect 509470 2790 509522 2796
rect 509988 1086 510016 2858
rect 510586 2802 510614 3060
rect 510540 2774 510614 2802
rect 511690 2802 511718 3060
rect 512794 2802 512822 3060
rect 513898 2802 513926 3060
rect 515002 2802 515030 3060
rect 516106 2802 516134 3060
rect 511690 2774 511764 2802
rect 512794 2774 512868 2802
rect 513898 2774 513972 2802
rect 515002 2774 515076 2802
rect 509976 1080 510028 1086
rect 509976 1022 510028 1028
rect 507860 1012 507912 1018
rect 507860 954 507912 960
rect 507308 876 507360 882
rect 507308 818 507360 824
rect 506480 740 506532 746
rect 506480 682 506532 688
rect 506112 536 506164 542
rect 505008 264 505060 270
rect 505008 206 505060 212
rect 505346 -960 505458 480
rect 506112 478 506164 484
rect 506492 480 506520 682
rect 506450 -960 506562 480
rect 507492 128 507544 134
rect 507646 82 507758 480
rect 507544 76 507758 82
rect 507492 70 507758 76
rect 507504 54 507758 70
rect 507646 -960 507758 54
rect 508842 218 508954 480
rect 509884 468 509936 474
rect 509884 410 509936 416
rect 509896 354 509924 410
rect 510038 354 510150 480
rect 509896 326 510150 354
rect 508842 202 509096 218
rect 508842 196 509108 202
rect 508842 190 509056 196
rect 508842 -960 508954 190
rect 509056 138 509108 144
rect 510038 -960 510150 326
rect 510540 134 510568 2774
rect 511264 672 511316 678
rect 511264 614 511316 620
rect 511276 480 511304 614
rect 510528 128 510580 134
rect 510528 70 510580 76
rect 511234 -960 511346 480
rect 511736 202 511764 2774
rect 512460 808 512512 814
rect 512460 750 512512 756
rect 512472 480 512500 750
rect 511724 196 511776 202
rect 511724 138 511776 144
rect 512430 -960 512542 480
rect 512840 474 512868 2774
rect 513944 678 513972 2774
rect 515048 746 515076 2774
rect 516060 2774 516134 2802
rect 517210 2802 517238 3060
rect 518314 2802 518342 3060
rect 519418 2802 519446 3060
rect 520522 2802 520550 3060
rect 521626 2802 521654 3060
rect 517210 2774 517284 2802
rect 518314 2774 518480 2802
rect 519418 2774 519492 2802
rect 520522 2774 520596 2802
rect 515036 740 515088 746
rect 515036 682 515088 688
rect 513932 672 513984 678
rect 513932 614 513984 620
rect 516060 626 516088 2774
rect 517256 814 517284 2774
rect 518256 944 518308 950
rect 518256 886 518308 892
rect 517244 808 517296 814
rect 517244 750 517296 756
rect 518268 626 518296 886
rect 516060 598 516180 626
rect 515772 536 515824 542
rect 512828 468 512880 474
rect 512828 410 512880 416
rect 513534 354 513646 480
rect 513392 338 513646 354
rect 513380 332 513646 338
rect 513432 326 513646 332
rect 513380 274 513432 280
rect 513534 -960 513646 326
rect 514730 354 514842 480
rect 515772 478 515824 484
rect 514944 400 514996 406
rect 514730 348 514944 354
rect 514730 342 514996 348
rect 515784 354 515812 478
rect 515926 354 516038 480
rect 516152 406 516180 598
rect 517152 604 517204 610
rect 518268 598 518388 626
rect 518452 610 518480 2774
rect 519464 678 519492 2774
rect 520568 1018 520596 2774
rect 521580 2774 521654 2802
rect 522730 2802 522758 3060
rect 523834 2922 523862 3060
rect 523822 2916 523874 2922
rect 523822 2858 523874 2864
rect 524938 2854 524966 3060
rect 525708 2916 525760 2922
rect 525708 2858 525760 2864
rect 524236 2848 524288 2854
rect 522730 2774 522804 2802
rect 524236 2790 524288 2796
rect 524926 2848 524978 2854
rect 524926 2790 524978 2796
rect 520556 1012 520608 1018
rect 520556 954 520608 960
rect 520740 944 520792 950
rect 520740 886 520792 892
rect 519452 672 519504 678
rect 519452 614 519504 620
rect 517152 546 517204 552
rect 517164 480 517192 546
rect 518360 480 518388 598
rect 518440 604 518492 610
rect 518440 546 518492 552
rect 520752 480 520780 886
rect 514730 326 514984 342
rect 515784 326 516038 354
rect 516140 400 516192 406
rect 516140 342 516192 348
rect 514730 -960 514842 326
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 218 519626 480
rect 519728 264 519780 270
rect 519514 212 519728 218
rect 519514 206 519780 212
rect 519514 190 519768 206
rect 519514 -960 519626 190
rect 520710 -960 520822 480
rect 521580 270 521608 2774
rect 521844 876 521896 882
rect 521844 818 521896 824
rect 521856 480 521884 818
rect 521568 264 521620 270
rect 521568 206 521620 212
rect 521814 -960 521926 480
rect 522776 338 522804 2774
rect 523040 1080 523092 1086
rect 523040 1022 523092 1028
rect 523052 480 523080 1022
rect 524248 480 524276 2790
rect 525720 1086 525748 2858
rect 526042 2802 526070 3060
rect 527146 2802 527174 3060
rect 526042 2774 526116 2802
rect 525708 1080 525760 1086
rect 525708 1022 525760 1028
rect 526088 950 526116 2774
rect 527100 2774 527174 2802
rect 528250 2802 528278 3060
rect 529354 2802 529382 3060
rect 530458 2802 530486 3060
rect 531562 2802 531590 3060
rect 532666 2802 532694 3060
rect 528250 2774 528324 2802
rect 529354 2774 529428 2802
rect 530458 2774 530532 2802
rect 531562 2774 531636 2802
rect 526076 944 526128 950
rect 526076 886 526128 892
rect 522764 332 522816 338
rect 522764 274 522816 280
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 82 525514 480
rect 526598 218 526710 480
rect 526456 202 526710 218
rect 526444 196 526710 202
rect 526496 190 526710 196
rect 526444 138 526496 144
rect 525616 128 525668 134
rect 525402 76 525616 82
rect 525402 70 525668 76
rect 525402 54 525656 70
rect 525402 -960 525514 54
rect 526598 -960 526710 190
rect 527100 134 527128 2774
rect 527794 354 527906 480
rect 528008 468 528060 474
rect 528008 410 528060 416
rect 528020 354 528048 410
rect 527794 326 528048 354
rect 527088 128 527140 134
rect 527088 70 527140 76
rect 527794 -960 527906 326
rect 528296 202 528324 2774
rect 529020 604 529072 610
rect 529020 546 529072 552
rect 529032 480 529060 546
rect 528284 196 528336 202
rect 528284 138 528336 144
rect 528990 -960 529102 480
rect 529400 474 529428 2774
rect 530504 746 530532 2774
rect 531608 882 531636 2774
rect 532620 2774 532694 2802
rect 533770 2802 533798 3060
rect 534874 2802 534902 3060
rect 535978 2802 536006 3060
rect 537082 2802 537110 3060
rect 538186 2802 538214 3060
rect 533770 2774 533936 2802
rect 534874 2774 535040 2802
rect 535978 2774 536052 2802
rect 537082 2774 537156 2802
rect 531596 876 531648 882
rect 531596 818 531648 824
rect 532332 808 532384 814
rect 532332 750 532384 756
rect 530124 740 530176 746
rect 530124 682 530176 688
rect 530492 740 530544 746
rect 530492 682 530544 688
rect 530136 480 530164 682
rect 529388 468 529440 474
rect 529388 410 529440 416
rect 530094 -960 530206 480
rect 531290 354 531402 480
rect 531504 400 531556 406
rect 531290 348 531504 354
rect 531290 342 531556 348
rect 532344 354 532372 750
rect 532620 746 532648 2774
rect 532608 740 532660 746
rect 532608 682 532660 688
rect 533712 604 533764 610
rect 533712 546 533764 552
rect 533724 480 533752 546
rect 532486 354 532598 480
rect 531290 326 531544 342
rect 532344 326 532598 354
rect 531290 -960 531402 326
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 533908 406 533936 2774
rect 534816 672 534868 678
rect 534868 620 534948 626
rect 534816 614 534948 620
rect 534828 598 534948 614
rect 535012 610 535040 2774
rect 536024 678 536052 2774
rect 537128 1222 537156 2774
rect 538140 2774 538214 2802
rect 539290 2802 539318 3060
rect 540394 2922 540422 3060
rect 541498 2922 541526 3060
rect 540382 2916 540434 2922
rect 540382 2858 540434 2864
rect 541348 2916 541400 2922
rect 541348 2858 541400 2864
rect 541486 2916 541538 2922
rect 541486 2858 541538 2864
rect 540796 2848 540848 2854
rect 539290 2774 539364 2802
rect 540796 2790 540848 2796
rect 537116 1216 537168 1222
rect 537116 1158 537168 1164
rect 536104 1012 536156 1018
rect 536104 954 536156 960
rect 536012 672 536064 678
rect 536012 614 536064 620
rect 534920 480 534948 598
rect 535000 604 535052 610
rect 535000 546 535052 552
rect 536116 480 536144 954
rect 533896 400 533948 406
rect 533896 342 533948 348
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 218 537290 480
rect 538140 270 538168 2774
rect 538374 354 538486 480
rect 538232 338 538486 354
rect 539336 338 539364 2774
rect 539600 1080 539652 1086
rect 539600 1022 539652 1028
rect 539612 480 539640 1022
rect 540808 480 540836 2790
rect 541360 1154 541388 2858
rect 542602 2802 542630 3060
rect 543706 2802 543734 3060
rect 542602 2774 542676 2802
rect 541348 1148 541400 1154
rect 541348 1090 541400 1096
rect 541992 944 542044 950
rect 541992 886 542044 892
rect 542004 480 542032 886
rect 542648 814 542676 2774
rect 543660 2774 543734 2802
rect 544810 2802 544838 3060
rect 545914 2802 545942 3060
rect 547018 2802 547046 3060
rect 548122 2802 548150 3060
rect 549226 2802 549254 3060
rect 544810 2774 544884 2802
rect 545914 2774 545988 2802
rect 547018 2774 547092 2802
rect 548122 2774 548196 2802
rect 542636 808 542688 814
rect 542636 750 542688 756
rect 538220 332 538486 338
rect 538272 326 538486 332
rect 538220 274 538272 280
rect 537392 264 537444 270
rect 537178 212 537392 218
rect 537178 206 537444 212
rect 538128 264 538180 270
rect 538128 206 538180 212
rect 537178 190 537432 206
rect 537178 -960 537290 190
rect 538374 -960 538486 326
rect 539324 332 539376 338
rect 539324 274 539376 280
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543004 128 543056 134
rect 543158 82 543270 480
rect 543660 134 543688 2774
rect 544354 218 544466 480
rect 544354 202 544608 218
rect 544856 202 544884 2774
rect 545960 950 545988 2774
rect 547064 1018 547092 2774
rect 548168 1086 548196 2774
rect 549180 2774 549254 2802
rect 550330 2802 550358 3060
rect 551434 2802 551462 3060
rect 550330 2774 550404 2802
rect 548156 1080 548208 1086
rect 548156 1022 548208 1028
rect 547052 1012 547104 1018
rect 547052 954 547104 960
rect 545948 944 546000 950
rect 545948 886 546000 892
rect 547880 876 547932 882
rect 547880 818 547932 824
rect 546684 740 546736 746
rect 546684 682 546736 688
rect 546696 480 546724 682
rect 547892 480 547920 818
rect 549180 626 549208 2774
rect 549076 604 549128 610
rect 549180 598 549300 626
rect 550376 610 550404 2774
rect 551388 2774 551462 2802
rect 552538 2802 552566 3060
rect 553642 2802 553670 3060
rect 554746 2802 554774 3060
rect 552538 2774 552612 2802
rect 551388 746 551416 2774
rect 552584 882 552612 2774
rect 553596 2774 553670 2802
rect 554608 2774 554774 2802
rect 555850 2802 555878 3060
rect 556436 2916 556488 2922
rect 556436 2858 556488 2864
rect 555850 2774 555924 2802
rect 552572 876 552624 882
rect 552572 818 552624 824
rect 551376 740 551428 746
rect 551376 682 551428 688
rect 551192 672 551244 678
rect 551244 620 551508 626
rect 551192 614 551508 620
rect 549076 546 549128 552
rect 549088 480 549116 546
rect 545458 354 545570 480
rect 545672 468 545724 474
rect 545672 410 545724 416
rect 545684 354 545712 410
rect 545458 326 545712 354
rect 544354 196 544620 202
rect 544354 190 544568 196
rect 543056 76 543270 82
rect 543004 70 543270 76
rect 543648 128 543700 134
rect 543648 70 543700 76
rect 543016 54 543270 70
rect 543158 -960 543270 54
rect 544354 -960 544466 190
rect 544568 138 544620 144
rect 544844 196 544896 202
rect 544844 138 544896 144
rect 545458 -960 545570 326
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 549272 406 549300 598
rect 550272 604 550324 610
rect 550272 546 550324 552
rect 550364 604 550416 610
rect 551204 598 551508 614
rect 550364 546 550416 552
rect 550284 480 550312 546
rect 551480 480 551508 598
rect 552664 604 552716 610
rect 552664 546 552716 552
rect 552676 480 552704 546
rect 549260 400 549312 406
rect 549260 342 549312 348
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553596 241 553624 2774
rect 553768 1216 553820 1222
rect 553768 1158 553820 1164
rect 553780 480 553808 1158
rect 553582 232 553638 241
rect 553582 167 553638 176
rect 553738 -960 553850 480
rect 554608 105 554636 2774
rect 554780 264 554832 270
rect 554934 218 555046 480
rect 555896 406 555924 2774
rect 555884 400 555936 406
rect 555884 342 555936 348
rect 556130 354 556242 480
rect 554832 212 555046 218
rect 554780 206 555046 212
rect 554792 190 555046 206
rect 554594 96 554650 105
rect 554594 31 554650 40
rect 554934 -960 555046 190
rect 556130 338 556384 354
rect 556448 338 556476 2858
rect 556954 2802 556982 3060
rect 558058 2802 558086 3060
rect 559162 2802 559190 3060
rect 560266 2802 560294 3060
rect 556954 2774 557028 2802
rect 558058 2774 558132 2802
rect 559162 2774 559236 2802
rect 557000 542 557028 2774
rect 557356 1148 557408 1154
rect 557356 1090 557408 1096
rect 556988 536 557040 542
rect 556988 478 557040 484
rect 557368 480 557396 1090
rect 558104 678 558132 2774
rect 559208 814 559236 2774
rect 560220 2774 560294 2802
rect 561370 2802 561398 3060
rect 562474 2802 562502 3060
rect 563578 2802 563606 3060
rect 561370 2774 561444 2802
rect 562474 2774 562548 2802
rect 563578 2774 563652 2802
rect 559104 808 559156 814
rect 559104 750 559156 756
rect 559196 808 559248 814
rect 559196 750 559248 756
rect 558092 672 558144 678
rect 558092 614 558144 620
rect 556130 332 556396 338
rect 556130 326 556344 332
rect 556130 -960 556242 326
rect 556344 274 556396 280
rect 556436 332 556488 338
rect 556436 274 556488 280
rect 557326 -960 557438 480
rect 558522 354 558634 480
rect 559116 354 559144 750
rect 559718 354 559830 480
rect 558522 338 558776 354
rect 558522 332 558788 338
rect 558522 326 558736 332
rect 558522 -960 558634 326
rect 559116 326 559830 354
rect 560220 338 560248 2774
rect 558736 274 558788 280
rect 559718 -960 559830 326
rect 560208 332 560260 338
rect 560208 274 560260 280
rect 560668 128 560720 134
rect 560822 82 560934 480
rect 561416 134 561444 2774
rect 562018 218 562130 480
rect 562018 202 562272 218
rect 562520 202 562548 2774
rect 563244 944 563296 950
rect 563244 886 563296 892
rect 563256 480 563284 886
rect 562018 196 562284 202
rect 562018 190 562232 196
rect 560720 76 560934 82
rect 560668 70 560934 76
rect 561404 128 561456 134
rect 561404 70 561456 76
rect 560680 54 560934 70
rect 560822 -960 560934 54
rect 562018 -960 562130 190
rect 562232 138 562284 144
rect 562508 196 562560 202
rect 562508 138 562560 144
rect 563214 -960 563326 480
rect 563624 270 563652 2774
rect 565636 1080 565688 1086
rect 565636 1022 565688 1028
rect 564440 1012 564492 1018
rect 564440 954 564492 960
rect 564452 480 564480 954
rect 565648 480 565676 1022
rect 570328 876 570380 882
rect 570328 818 570380 824
rect 569132 740 569184 746
rect 569132 682 569184 688
rect 568028 604 568080 610
rect 568028 546 568080 552
rect 568040 480 568068 546
rect 569144 480 569172 682
rect 570340 480 570368 818
rect 577412 808 577464 814
rect 577412 750 577464 756
rect 576308 672 576360 678
rect 576308 614 576360 620
rect 575112 604 575164 610
rect 575112 546 575164 552
rect 575124 480 575152 546
rect 576320 480 576348 614
rect 577424 480 577452 750
rect 563612 264 563664 270
rect 563612 206 563664 212
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 354 566914 480
rect 567016 468 567068 474
rect 567016 410 567068 416
rect 567028 354 567056 410
rect 566802 326 567056 354
rect 566802 -960 566914 326
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571338 232 571394 241
rect 571494 218 571606 480
rect 571394 190 571606 218
rect 571338 167 571394 176
rect 571494 -960 571606 190
rect 572690 82 572802 480
rect 573732 400 573784 406
rect 573886 354 573998 480
rect 573784 348 573998 354
rect 573732 342 573998 348
rect 573744 326 573998 342
rect 572902 96 572958 105
rect 572690 54 572902 82
rect 572690 -960 572802 54
rect 572902 31 572958 40
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 354 578690 480
rect 578578 338 578832 354
rect 578578 332 578844 338
rect 578578 326 578792 332
rect 578578 -960 578690 326
rect 578792 274 578844 280
rect 579774 -960 579886 480
rect 580970 82 581082 480
rect 582166 218 582278 480
rect 582024 202 582278 218
rect 582012 196 582278 202
rect 582064 190 582278 196
rect 582012 138 582064 144
rect 581184 128 581236 134
rect 580970 76 581184 82
rect 580970 70 581236 76
rect 580970 54 581224 70
rect 580970 -960 581082 54
rect 582166 -960 582278 190
rect 583362 218 583474 480
rect 583576 264 583628 270
rect 583362 212 583576 218
rect 583362 206 583628 212
rect 583362 190 583616 206
rect 583362 -960 583474 190
<< via2 >>
rect 3882 448 3938 504
rect 16210 40 16266 96
rect 20442 312 20498 368
rect 22006 176 22062 232
rect 23662 448 23718 504
rect 34426 40 34482 96
rect 39118 312 39174 368
rect 39394 40 39450 96
rect 40222 176 40278 232
rect 45282 176 45338 232
rect 56782 40 56838 96
rect 62394 176 62450 232
rect 553582 176 553638 232
rect 554594 40 554650 96
rect 571338 176 571394 232
rect 572902 40 572958 96
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
rect 3877 506 3943 509
rect 23657 506 23723 509
rect 3877 504 23723 506
rect 3877 448 3882 504
rect 3938 448 23662 504
rect 23718 448 23723 504
rect 3877 446 23723 448
rect 3877 443 3943 446
rect 23657 443 23723 446
rect 20437 370 20503 373
rect 39113 370 39179 373
rect 20437 368 39179 370
rect 20437 312 20442 368
rect 20498 312 39118 368
rect 39174 312 39179 368
rect 20437 310 39179 312
rect 20437 307 20503 310
rect 39113 307 39179 310
rect 22001 234 22067 237
rect 40217 234 40283 237
rect 22001 232 40283 234
rect 22001 176 22006 232
rect 22062 176 40222 232
rect 40278 176 40283 232
rect 22001 174 40283 176
rect 22001 171 22067 174
rect 40217 171 40283 174
rect 45277 234 45343 237
rect 62389 234 62455 237
rect 45277 232 62455 234
rect 45277 176 45282 232
rect 45338 176 62394 232
rect 62450 176 62455 232
rect 45277 174 62455 176
rect 45277 171 45343 174
rect 62389 171 62455 174
rect 553577 234 553643 237
rect 571333 234 571399 237
rect 553577 232 571399 234
rect 553577 176 553582 232
rect 553638 176 571338 232
rect 571394 176 571399 232
rect 553577 174 571399 176
rect 553577 171 553643 174
rect 571333 171 571399 174
rect 16205 98 16271 101
rect 34421 98 34487 101
rect 16205 96 34487 98
rect 16205 40 16210 96
rect 16266 40 34426 96
rect 34482 40 34487 96
rect 16205 38 34487 40
rect 16205 35 16271 38
rect 34421 35 34487 38
rect 39389 98 39455 101
rect 56777 98 56843 101
rect 39389 96 56843 98
rect 39389 40 39394 96
rect 39450 40 56782 96
rect 56838 40 56843 96
rect 39389 38 56843 40
rect 39389 35 39455 38
rect 56777 35 56843 38
rect 554589 98 554655 101
rect 572897 98 572963 101
rect 554589 96 572963 98
rect 554589 40 554594 96
rect 554650 40 572902 96
rect 572958 40 572963 96
rect 554589 38 572963 40
rect 554589 35 554655 38
rect 572897 35 572963 38
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711002 -8694 711558
rect -8138 711002 -8106 711558
rect -8726 677494 -8106 711002
rect -8726 676938 -8694 677494
rect -8138 676938 -8106 677494
rect -8726 641494 -8106 676938
rect -8726 640938 -8694 641494
rect -8138 640938 -8106 641494
rect -8726 605494 -8106 640938
rect -8726 604938 -8694 605494
rect -8138 604938 -8106 605494
rect -8726 569494 -8106 604938
rect -8726 568938 -8694 569494
rect -8138 568938 -8106 569494
rect -8726 533494 -8106 568938
rect -8726 532938 -8694 533494
rect -8138 532938 -8106 533494
rect -8726 497494 -8106 532938
rect -8726 496938 -8694 497494
rect -8138 496938 -8106 497494
rect -8726 461494 -8106 496938
rect -8726 460938 -8694 461494
rect -8138 460938 -8106 461494
rect -8726 425494 -8106 460938
rect -8726 424938 -8694 425494
rect -8138 424938 -8106 425494
rect -8726 389494 -8106 424938
rect -8726 388938 -8694 389494
rect -8138 388938 -8106 389494
rect -8726 353494 -8106 388938
rect -8726 352938 -8694 353494
rect -8138 352938 -8106 353494
rect -8726 317494 -8106 352938
rect -8726 316938 -8694 317494
rect -8138 316938 -8106 317494
rect -8726 281494 -8106 316938
rect -8726 280938 -8694 281494
rect -8138 280938 -8106 281494
rect -8726 245494 -8106 280938
rect -8726 244938 -8694 245494
rect -8138 244938 -8106 245494
rect -8726 209494 -8106 244938
rect -8726 208938 -8694 209494
rect -8138 208938 -8106 209494
rect -8726 173494 -8106 208938
rect -8726 172938 -8694 173494
rect -8138 172938 -8106 173494
rect -8726 137494 -8106 172938
rect -8726 136938 -8694 137494
rect -8138 136938 -8106 137494
rect -8726 101494 -8106 136938
rect -8726 100938 -8694 101494
rect -8138 100938 -8106 101494
rect -8726 65494 -8106 100938
rect -8726 64938 -8694 65494
rect -8138 64938 -8106 65494
rect -8726 29494 -8106 64938
rect -8726 28938 -8694 29494
rect -8138 28938 -8106 29494
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710042 -7734 710598
rect -7178 710042 -7146 710598
rect -7766 673774 -7146 710042
rect -7766 673218 -7734 673774
rect -7178 673218 -7146 673774
rect -7766 637774 -7146 673218
rect -7766 637218 -7734 637774
rect -7178 637218 -7146 637774
rect -7766 601774 -7146 637218
rect -7766 601218 -7734 601774
rect -7178 601218 -7146 601774
rect -7766 565774 -7146 601218
rect -7766 565218 -7734 565774
rect -7178 565218 -7146 565774
rect -7766 529774 -7146 565218
rect -7766 529218 -7734 529774
rect -7178 529218 -7146 529774
rect -7766 493774 -7146 529218
rect -7766 493218 -7734 493774
rect -7178 493218 -7146 493774
rect -7766 457774 -7146 493218
rect -7766 457218 -7734 457774
rect -7178 457218 -7146 457774
rect -7766 421774 -7146 457218
rect -7766 421218 -7734 421774
rect -7178 421218 -7146 421774
rect -7766 385774 -7146 421218
rect -7766 385218 -7734 385774
rect -7178 385218 -7146 385774
rect -7766 349774 -7146 385218
rect -7766 349218 -7734 349774
rect -7178 349218 -7146 349774
rect -7766 313774 -7146 349218
rect -7766 313218 -7734 313774
rect -7178 313218 -7146 313774
rect -7766 277774 -7146 313218
rect -7766 277218 -7734 277774
rect -7178 277218 -7146 277774
rect -7766 241774 -7146 277218
rect -7766 241218 -7734 241774
rect -7178 241218 -7146 241774
rect -7766 205774 -7146 241218
rect -7766 205218 -7734 205774
rect -7178 205218 -7146 205774
rect -7766 169774 -7146 205218
rect -7766 169218 -7734 169774
rect -7178 169218 -7146 169774
rect -7766 133774 -7146 169218
rect -7766 133218 -7734 133774
rect -7178 133218 -7146 133774
rect -7766 97774 -7146 133218
rect -7766 97218 -7734 97774
rect -7178 97218 -7146 97774
rect -7766 61774 -7146 97218
rect -7766 61218 -7734 61774
rect -7178 61218 -7146 61774
rect -7766 25774 -7146 61218
rect -7766 25218 -7734 25774
rect -7178 25218 -7146 25774
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709082 -6774 709638
rect -6218 709082 -6186 709638
rect -6806 670054 -6186 709082
rect -6806 669498 -6774 670054
rect -6218 669498 -6186 670054
rect -6806 634054 -6186 669498
rect -6806 633498 -6774 634054
rect -6218 633498 -6186 634054
rect -6806 598054 -6186 633498
rect -6806 597498 -6774 598054
rect -6218 597498 -6186 598054
rect -6806 562054 -6186 597498
rect -6806 561498 -6774 562054
rect -6218 561498 -6186 562054
rect -6806 526054 -6186 561498
rect -6806 525498 -6774 526054
rect -6218 525498 -6186 526054
rect -6806 490054 -6186 525498
rect -6806 489498 -6774 490054
rect -6218 489498 -6186 490054
rect -6806 454054 -6186 489498
rect -6806 453498 -6774 454054
rect -6218 453498 -6186 454054
rect -6806 418054 -6186 453498
rect -6806 417498 -6774 418054
rect -6218 417498 -6186 418054
rect -6806 382054 -6186 417498
rect -6806 381498 -6774 382054
rect -6218 381498 -6186 382054
rect -6806 346054 -6186 381498
rect -6806 345498 -6774 346054
rect -6218 345498 -6186 346054
rect -6806 310054 -6186 345498
rect -6806 309498 -6774 310054
rect -6218 309498 -6186 310054
rect -6806 274054 -6186 309498
rect -6806 273498 -6774 274054
rect -6218 273498 -6186 274054
rect -6806 238054 -6186 273498
rect -6806 237498 -6774 238054
rect -6218 237498 -6186 238054
rect -6806 202054 -6186 237498
rect -6806 201498 -6774 202054
rect -6218 201498 -6186 202054
rect -6806 166054 -6186 201498
rect -6806 165498 -6774 166054
rect -6218 165498 -6186 166054
rect -6806 130054 -6186 165498
rect -6806 129498 -6774 130054
rect -6218 129498 -6186 130054
rect -6806 94054 -6186 129498
rect -6806 93498 -6774 94054
rect -6218 93498 -6186 94054
rect -6806 58054 -6186 93498
rect -6806 57498 -6774 58054
rect -6218 57498 -6186 58054
rect -6806 22054 -6186 57498
rect -6806 21498 -6774 22054
rect -6218 21498 -6186 22054
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708122 -5814 708678
rect -5258 708122 -5226 708678
rect -5846 666334 -5226 708122
rect -5846 665778 -5814 666334
rect -5258 665778 -5226 666334
rect -5846 630334 -5226 665778
rect -5846 629778 -5814 630334
rect -5258 629778 -5226 630334
rect -5846 594334 -5226 629778
rect -5846 593778 -5814 594334
rect -5258 593778 -5226 594334
rect -5846 558334 -5226 593778
rect -5846 557778 -5814 558334
rect -5258 557778 -5226 558334
rect -5846 522334 -5226 557778
rect -5846 521778 -5814 522334
rect -5258 521778 -5226 522334
rect -5846 486334 -5226 521778
rect -5846 485778 -5814 486334
rect -5258 485778 -5226 486334
rect -5846 450334 -5226 485778
rect -5846 449778 -5814 450334
rect -5258 449778 -5226 450334
rect -5846 414334 -5226 449778
rect -5846 413778 -5814 414334
rect -5258 413778 -5226 414334
rect -5846 378334 -5226 413778
rect -5846 377778 -5814 378334
rect -5258 377778 -5226 378334
rect -5846 342334 -5226 377778
rect -5846 341778 -5814 342334
rect -5258 341778 -5226 342334
rect -5846 306334 -5226 341778
rect -5846 305778 -5814 306334
rect -5258 305778 -5226 306334
rect -5846 270334 -5226 305778
rect -5846 269778 -5814 270334
rect -5258 269778 -5226 270334
rect -5846 234334 -5226 269778
rect -5846 233778 -5814 234334
rect -5258 233778 -5226 234334
rect -5846 198334 -5226 233778
rect -5846 197778 -5814 198334
rect -5258 197778 -5226 198334
rect -5846 162334 -5226 197778
rect -5846 161778 -5814 162334
rect -5258 161778 -5226 162334
rect -5846 126334 -5226 161778
rect -5846 125778 -5814 126334
rect -5258 125778 -5226 126334
rect -5846 90334 -5226 125778
rect -5846 89778 -5814 90334
rect -5258 89778 -5226 90334
rect -5846 54334 -5226 89778
rect -5846 53778 -5814 54334
rect -5258 53778 -5226 54334
rect -5846 18334 -5226 53778
rect -5846 17778 -5814 18334
rect -5258 17778 -5226 18334
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707162 -4854 707718
rect -4298 707162 -4266 707718
rect -4886 698614 -4266 707162
rect -4886 698058 -4854 698614
rect -4298 698058 -4266 698614
rect -4886 662614 -4266 698058
rect -4886 662058 -4854 662614
rect -4298 662058 -4266 662614
rect -4886 626614 -4266 662058
rect -4886 626058 -4854 626614
rect -4298 626058 -4266 626614
rect -4886 590614 -4266 626058
rect -4886 590058 -4854 590614
rect -4298 590058 -4266 590614
rect -4886 554614 -4266 590058
rect -4886 554058 -4854 554614
rect -4298 554058 -4266 554614
rect -4886 518614 -4266 554058
rect -4886 518058 -4854 518614
rect -4298 518058 -4266 518614
rect -4886 482614 -4266 518058
rect -4886 482058 -4854 482614
rect -4298 482058 -4266 482614
rect -4886 446614 -4266 482058
rect -4886 446058 -4854 446614
rect -4298 446058 -4266 446614
rect -4886 410614 -4266 446058
rect -4886 410058 -4854 410614
rect -4298 410058 -4266 410614
rect -4886 374614 -4266 410058
rect -4886 374058 -4854 374614
rect -4298 374058 -4266 374614
rect -4886 338614 -4266 374058
rect -4886 338058 -4854 338614
rect -4298 338058 -4266 338614
rect -4886 302614 -4266 338058
rect -4886 302058 -4854 302614
rect -4298 302058 -4266 302614
rect -4886 266614 -4266 302058
rect -4886 266058 -4854 266614
rect -4298 266058 -4266 266614
rect -4886 230614 -4266 266058
rect -4886 230058 -4854 230614
rect -4298 230058 -4266 230614
rect -4886 194614 -4266 230058
rect -4886 194058 -4854 194614
rect -4298 194058 -4266 194614
rect -4886 158614 -4266 194058
rect -4886 158058 -4854 158614
rect -4298 158058 -4266 158614
rect -4886 122614 -4266 158058
rect -4886 122058 -4854 122614
rect -4298 122058 -4266 122614
rect -4886 86614 -4266 122058
rect -4886 86058 -4854 86614
rect -4298 86058 -4266 86614
rect -4886 50614 -4266 86058
rect -4886 50058 -4854 50614
rect -4298 50058 -4266 50614
rect -4886 14614 -4266 50058
rect -4886 14058 -4854 14614
rect -4298 14058 -4266 14614
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706202 -3894 706758
rect -3338 706202 -3306 706758
rect -3926 694894 -3306 706202
rect -3926 694338 -3894 694894
rect -3338 694338 -3306 694894
rect -3926 658894 -3306 694338
rect -3926 658338 -3894 658894
rect -3338 658338 -3306 658894
rect -3926 622894 -3306 658338
rect -3926 622338 -3894 622894
rect -3338 622338 -3306 622894
rect -3926 586894 -3306 622338
rect -3926 586338 -3894 586894
rect -3338 586338 -3306 586894
rect -3926 550894 -3306 586338
rect -3926 550338 -3894 550894
rect -3338 550338 -3306 550894
rect -3926 514894 -3306 550338
rect -3926 514338 -3894 514894
rect -3338 514338 -3306 514894
rect -3926 478894 -3306 514338
rect -3926 478338 -3894 478894
rect -3338 478338 -3306 478894
rect -3926 442894 -3306 478338
rect -3926 442338 -3894 442894
rect -3338 442338 -3306 442894
rect -3926 406894 -3306 442338
rect -3926 406338 -3894 406894
rect -3338 406338 -3306 406894
rect -3926 370894 -3306 406338
rect -3926 370338 -3894 370894
rect -3338 370338 -3306 370894
rect -3926 334894 -3306 370338
rect -3926 334338 -3894 334894
rect -3338 334338 -3306 334894
rect -3926 298894 -3306 334338
rect -3926 298338 -3894 298894
rect -3338 298338 -3306 298894
rect -3926 262894 -3306 298338
rect -3926 262338 -3894 262894
rect -3338 262338 -3306 262894
rect -3926 226894 -3306 262338
rect -3926 226338 -3894 226894
rect -3338 226338 -3306 226894
rect -3926 190894 -3306 226338
rect -3926 190338 -3894 190894
rect -3338 190338 -3306 190894
rect -3926 154894 -3306 190338
rect -3926 154338 -3894 154894
rect -3338 154338 -3306 154894
rect -3926 118894 -3306 154338
rect -3926 118338 -3894 118894
rect -3338 118338 -3306 118894
rect -3926 82894 -3306 118338
rect -3926 82338 -3894 82894
rect -3338 82338 -3306 82894
rect -3926 46894 -3306 82338
rect -3926 46338 -3894 46894
rect -3338 46338 -3306 46894
rect -3926 10894 -3306 46338
rect -3926 10338 -3894 10894
rect -3338 10338 -3306 10894
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705242 -2934 705798
rect -2378 705242 -2346 705798
rect -2966 691174 -2346 705242
rect -2966 690618 -2934 691174
rect -2378 690618 -2346 691174
rect -2966 655174 -2346 690618
rect -2966 654618 -2934 655174
rect -2378 654618 -2346 655174
rect -2966 619174 -2346 654618
rect -2966 618618 -2934 619174
rect -2378 618618 -2346 619174
rect -2966 583174 -2346 618618
rect -2966 582618 -2934 583174
rect -2378 582618 -2346 583174
rect -2966 547174 -2346 582618
rect -2966 546618 -2934 547174
rect -2378 546618 -2346 547174
rect -2966 511174 -2346 546618
rect -2966 510618 -2934 511174
rect -2378 510618 -2346 511174
rect -2966 475174 -2346 510618
rect -2966 474618 -2934 475174
rect -2378 474618 -2346 475174
rect -2966 439174 -2346 474618
rect -2966 438618 -2934 439174
rect -2378 438618 -2346 439174
rect -2966 403174 -2346 438618
rect -2966 402618 -2934 403174
rect -2378 402618 -2346 403174
rect -2966 367174 -2346 402618
rect -2966 366618 -2934 367174
rect -2378 366618 -2346 367174
rect -2966 331174 -2346 366618
rect -2966 330618 -2934 331174
rect -2378 330618 -2346 331174
rect -2966 295174 -2346 330618
rect -2966 294618 -2934 295174
rect -2378 294618 -2346 295174
rect -2966 259174 -2346 294618
rect -2966 258618 -2934 259174
rect -2378 258618 -2346 259174
rect -2966 223174 -2346 258618
rect -2966 222618 -2934 223174
rect -2378 222618 -2346 223174
rect -2966 187174 -2346 222618
rect -2966 186618 -2934 187174
rect -2378 186618 -2346 187174
rect -2966 151174 -2346 186618
rect -2966 150618 -2934 151174
rect -2378 150618 -2346 151174
rect -2966 115174 -2346 150618
rect -2966 114618 -2934 115174
rect -2378 114618 -2346 115174
rect -2966 79174 -2346 114618
rect -2966 78618 -2934 79174
rect -2378 78618 -2346 79174
rect -2966 43174 -2346 78618
rect -2966 42618 -2934 43174
rect -2378 42618 -2346 43174
rect -2966 7174 -2346 42618
rect -2966 6618 -2934 7174
rect -2378 6618 -2346 7174
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704282 -1974 704838
rect -1418 704282 -1386 704838
rect -2006 687454 -1386 704282
rect -2006 686898 -1974 687454
rect -1418 686898 -1386 687454
rect -2006 651454 -1386 686898
rect -2006 650898 -1974 651454
rect -1418 650898 -1386 651454
rect -2006 615454 -1386 650898
rect -2006 614898 -1974 615454
rect -1418 614898 -1386 615454
rect -2006 579454 -1386 614898
rect -2006 578898 -1974 579454
rect -1418 578898 -1386 579454
rect -2006 543454 -1386 578898
rect -2006 542898 -1974 543454
rect -1418 542898 -1386 543454
rect -2006 507454 -1386 542898
rect -2006 506898 -1974 507454
rect -1418 506898 -1386 507454
rect -2006 471454 -1386 506898
rect -2006 470898 -1974 471454
rect -1418 470898 -1386 471454
rect -2006 435454 -1386 470898
rect -2006 434898 -1974 435454
rect -1418 434898 -1386 435454
rect -2006 399454 -1386 434898
rect -2006 398898 -1974 399454
rect -1418 398898 -1386 399454
rect -2006 363454 -1386 398898
rect -2006 362898 -1974 363454
rect -1418 362898 -1386 363454
rect -2006 327454 -1386 362898
rect -2006 326898 -1974 327454
rect -1418 326898 -1386 327454
rect -2006 291454 -1386 326898
rect -2006 290898 -1974 291454
rect -1418 290898 -1386 291454
rect -2006 255454 -1386 290898
rect -2006 254898 -1974 255454
rect -1418 254898 -1386 255454
rect -2006 219454 -1386 254898
rect -2006 218898 -1974 219454
rect -1418 218898 -1386 219454
rect -2006 183454 -1386 218898
rect -2006 182898 -1974 183454
rect -1418 182898 -1386 183454
rect -2006 147454 -1386 182898
rect -2006 146898 -1974 147454
rect -1418 146898 -1386 147454
rect -2006 111454 -1386 146898
rect -2006 110898 -1974 111454
rect -1418 110898 -1386 111454
rect -2006 75454 -1386 110898
rect -2006 74898 -1974 75454
rect -1418 74898 -1386 75454
rect -2006 39454 -1386 74898
rect -2006 38898 -1974 39454
rect -1418 38898 -1386 39454
rect -2006 3454 -1386 38898
rect -2006 2898 -1974 3454
rect -1418 2898 -1386 3454
rect -2006 -346 -1386 2898
rect -2006 -902 -1974 -346
rect -1418 -902 -1386 -346
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704282 1826 704838
rect 2382 704282 2414 704838
rect 1794 687454 2414 704282
rect 1794 686898 1826 687454
rect 2382 686898 2414 687454
rect 1794 651454 2414 686898
rect 1794 650898 1826 651454
rect 2382 650898 2414 651454
rect 1794 615454 2414 650898
rect 1794 614898 1826 615454
rect 2382 614898 2414 615454
rect 1794 579454 2414 614898
rect 1794 578898 1826 579454
rect 2382 578898 2414 579454
rect 1794 543454 2414 578898
rect 1794 542898 1826 543454
rect 2382 542898 2414 543454
rect 1794 507454 2414 542898
rect 1794 506898 1826 507454
rect 2382 506898 2414 507454
rect 1794 471454 2414 506898
rect 1794 470898 1826 471454
rect 2382 470898 2414 471454
rect 1794 435454 2414 470898
rect 1794 434898 1826 435454
rect 2382 434898 2414 435454
rect 1794 399454 2414 434898
rect 1794 398898 1826 399454
rect 2382 398898 2414 399454
rect 1794 363454 2414 398898
rect 1794 362898 1826 363454
rect 2382 362898 2414 363454
rect 1794 327454 2414 362898
rect 1794 326898 1826 327454
rect 2382 326898 2414 327454
rect 1794 291454 2414 326898
rect 1794 290898 1826 291454
rect 2382 290898 2414 291454
rect 1794 255454 2414 290898
rect 1794 254898 1826 255454
rect 2382 254898 2414 255454
rect 1794 219454 2414 254898
rect 1794 218898 1826 219454
rect 2382 218898 2414 219454
rect 1794 183454 2414 218898
rect 1794 182898 1826 183454
rect 2382 182898 2414 183454
rect 1794 147454 2414 182898
rect 1794 146898 1826 147454
rect 2382 146898 2414 147454
rect 1794 111454 2414 146898
rect 1794 110898 1826 111454
rect 2382 110898 2414 111454
rect 1794 75454 2414 110898
rect 1794 74898 1826 75454
rect 2382 74898 2414 75454
rect 1794 39454 2414 74898
rect 1794 38898 1826 39454
rect 2382 38898 2414 39454
rect 1794 3454 2414 38898
rect 1794 2898 1826 3454
rect 2382 2898 2414 3454
rect 1794 -346 2414 2898
rect 1794 -902 1826 -346
rect 2382 -902 2414 -346
rect -2966 -1862 -2934 -1306
rect -2378 -1862 -2346 -1306
rect -2966 -1894 -2346 -1862
rect -3926 -2822 -3894 -2266
rect -3338 -2822 -3306 -2266
rect -3926 -2854 -3306 -2822
rect -4886 -3782 -4854 -3226
rect -4298 -3782 -4266 -3226
rect -4886 -3814 -4266 -3782
rect -5846 -4742 -5814 -4186
rect -5258 -4742 -5226 -4186
rect -5846 -4774 -5226 -4742
rect -6806 -5702 -6774 -5146
rect -6218 -5702 -6186 -5146
rect -6806 -5734 -6186 -5702
rect -7766 -6662 -7734 -6106
rect -7178 -6662 -7146 -6106
rect -7766 -6694 -7146 -6662
rect -8726 -7622 -8694 -7066
rect -8138 -7622 -8106 -7066
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 705798 6134 711590
rect 5514 705242 5546 705798
rect 6102 705242 6134 705798
rect 5514 691174 6134 705242
rect 5514 690618 5546 691174
rect 6102 690618 6134 691174
rect 5514 655174 6134 690618
rect 5514 654618 5546 655174
rect 6102 654618 6134 655174
rect 5514 619174 6134 654618
rect 5514 618618 5546 619174
rect 6102 618618 6134 619174
rect 5514 583174 6134 618618
rect 5514 582618 5546 583174
rect 6102 582618 6134 583174
rect 5514 547174 6134 582618
rect 5514 546618 5546 547174
rect 6102 546618 6134 547174
rect 5514 511174 6134 546618
rect 5514 510618 5546 511174
rect 6102 510618 6134 511174
rect 5514 475174 6134 510618
rect 5514 474618 5546 475174
rect 6102 474618 6134 475174
rect 5514 439174 6134 474618
rect 5514 438618 5546 439174
rect 6102 438618 6134 439174
rect 5514 403174 6134 438618
rect 5514 402618 5546 403174
rect 6102 402618 6134 403174
rect 5514 367174 6134 402618
rect 5514 366618 5546 367174
rect 6102 366618 6134 367174
rect 5514 331174 6134 366618
rect 5514 330618 5546 331174
rect 6102 330618 6134 331174
rect 5514 295174 6134 330618
rect 5514 294618 5546 295174
rect 6102 294618 6134 295174
rect 5514 259174 6134 294618
rect 5514 258618 5546 259174
rect 6102 258618 6134 259174
rect 5514 223174 6134 258618
rect 5514 222618 5546 223174
rect 6102 222618 6134 223174
rect 5514 187174 6134 222618
rect 5514 186618 5546 187174
rect 6102 186618 6134 187174
rect 5514 151174 6134 186618
rect 5514 150618 5546 151174
rect 6102 150618 6134 151174
rect 5514 115174 6134 150618
rect 5514 114618 5546 115174
rect 6102 114618 6134 115174
rect 5514 79174 6134 114618
rect 5514 78618 5546 79174
rect 6102 78618 6134 79174
rect 5514 43174 6134 78618
rect 5514 42618 5546 43174
rect 6102 42618 6134 43174
rect 5514 7174 6134 42618
rect 5514 6618 5546 7174
rect 6102 6618 6134 7174
rect 5514 -1306 6134 6618
rect 5514 -1862 5546 -1306
rect 6102 -1862 6134 -1306
rect 5514 -7654 6134 -1862
rect 9234 706758 9854 711590
rect 9234 706202 9266 706758
rect 9822 706202 9854 706758
rect 9234 694894 9854 706202
rect 9234 694338 9266 694894
rect 9822 694338 9854 694894
rect 9234 658894 9854 694338
rect 9234 658338 9266 658894
rect 9822 658338 9854 658894
rect 9234 622894 9854 658338
rect 9234 622338 9266 622894
rect 9822 622338 9854 622894
rect 9234 586894 9854 622338
rect 9234 586338 9266 586894
rect 9822 586338 9854 586894
rect 9234 550894 9854 586338
rect 9234 550338 9266 550894
rect 9822 550338 9854 550894
rect 9234 514894 9854 550338
rect 9234 514338 9266 514894
rect 9822 514338 9854 514894
rect 9234 478894 9854 514338
rect 9234 478338 9266 478894
rect 9822 478338 9854 478894
rect 9234 442894 9854 478338
rect 9234 442338 9266 442894
rect 9822 442338 9854 442894
rect 9234 406894 9854 442338
rect 9234 406338 9266 406894
rect 9822 406338 9854 406894
rect 9234 370894 9854 406338
rect 9234 370338 9266 370894
rect 9822 370338 9854 370894
rect 9234 334894 9854 370338
rect 9234 334338 9266 334894
rect 9822 334338 9854 334894
rect 9234 298894 9854 334338
rect 9234 298338 9266 298894
rect 9822 298338 9854 298894
rect 9234 262894 9854 298338
rect 9234 262338 9266 262894
rect 9822 262338 9854 262894
rect 9234 226894 9854 262338
rect 9234 226338 9266 226894
rect 9822 226338 9854 226894
rect 9234 190894 9854 226338
rect 9234 190338 9266 190894
rect 9822 190338 9854 190894
rect 9234 154894 9854 190338
rect 9234 154338 9266 154894
rect 9822 154338 9854 154894
rect 9234 118894 9854 154338
rect 9234 118338 9266 118894
rect 9822 118338 9854 118894
rect 9234 82894 9854 118338
rect 9234 82338 9266 82894
rect 9822 82338 9854 82894
rect 9234 46894 9854 82338
rect 9234 46338 9266 46894
rect 9822 46338 9854 46894
rect 9234 10894 9854 46338
rect 9234 10338 9266 10894
rect 9822 10338 9854 10894
rect 9234 -2266 9854 10338
rect 9234 -2822 9266 -2266
rect 9822 -2822 9854 -2266
rect 9234 -7654 9854 -2822
rect 12954 707718 13574 711590
rect 12954 707162 12986 707718
rect 13542 707162 13574 707718
rect 12954 698614 13574 707162
rect 12954 698058 12986 698614
rect 13542 698058 13574 698614
rect 12954 662614 13574 698058
rect 12954 662058 12986 662614
rect 13542 662058 13574 662614
rect 12954 626614 13574 662058
rect 12954 626058 12986 626614
rect 13542 626058 13574 626614
rect 12954 590614 13574 626058
rect 12954 590058 12986 590614
rect 13542 590058 13574 590614
rect 12954 554614 13574 590058
rect 12954 554058 12986 554614
rect 13542 554058 13574 554614
rect 12954 518614 13574 554058
rect 12954 518058 12986 518614
rect 13542 518058 13574 518614
rect 12954 482614 13574 518058
rect 12954 482058 12986 482614
rect 13542 482058 13574 482614
rect 12954 446614 13574 482058
rect 12954 446058 12986 446614
rect 13542 446058 13574 446614
rect 12954 410614 13574 446058
rect 12954 410058 12986 410614
rect 13542 410058 13574 410614
rect 12954 374614 13574 410058
rect 12954 374058 12986 374614
rect 13542 374058 13574 374614
rect 12954 338614 13574 374058
rect 12954 338058 12986 338614
rect 13542 338058 13574 338614
rect 12954 302614 13574 338058
rect 16674 708678 17294 711590
rect 16674 708122 16706 708678
rect 17262 708122 17294 708678
rect 16674 666334 17294 708122
rect 16674 665778 16706 666334
rect 17262 665778 17294 666334
rect 16674 630334 17294 665778
rect 16674 629778 16706 630334
rect 17262 629778 17294 630334
rect 16674 594334 17294 629778
rect 16674 593778 16706 594334
rect 17262 593778 17294 594334
rect 16674 558334 17294 593778
rect 16674 557778 16706 558334
rect 17262 557778 17294 558334
rect 16674 522334 17294 557778
rect 16674 521778 16706 522334
rect 17262 521778 17294 522334
rect 16674 486334 17294 521778
rect 16674 485778 16706 486334
rect 17262 485778 17294 486334
rect 16674 450334 17294 485778
rect 16674 449778 16706 450334
rect 17262 449778 17294 450334
rect 16674 414334 17294 449778
rect 16674 413778 16706 414334
rect 17262 413778 17294 414334
rect 16674 378334 17294 413778
rect 16674 377778 16706 378334
rect 17262 377778 17294 378334
rect 16674 342334 17294 377778
rect 16674 341778 16706 342334
rect 17262 341778 17294 342334
rect 16208 327454 16528 327486
rect 16208 327218 16250 327454
rect 16486 327218 16528 327454
rect 16208 327134 16528 327218
rect 16208 326898 16250 327134
rect 16486 326898 16528 327134
rect 16208 326866 16528 326898
rect 12954 302058 12986 302614
rect 13542 302058 13574 302614
rect 12954 266614 13574 302058
rect 16674 306334 17294 341778
rect 16674 305778 16706 306334
rect 17262 305778 17294 306334
rect 16208 291454 16528 291486
rect 16208 291218 16250 291454
rect 16486 291218 16528 291454
rect 16208 291134 16528 291218
rect 16208 290898 16250 291134
rect 16486 290898 16528 291134
rect 16208 290866 16528 290898
rect 12954 266058 12986 266614
rect 13542 266058 13574 266614
rect 12954 230614 13574 266058
rect 16674 270334 17294 305778
rect 16674 269778 16706 270334
rect 17262 269778 17294 270334
rect 16208 255454 16528 255486
rect 16208 255218 16250 255454
rect 16486 255218 16528 255454
rect 16208 255134 16528 255218
rect 16208 254898 16250 255134
rect 16486 254898 16528 255134
rect 16208 254866 16528 254898
rect 12954 230058 12986 230614
rect 13542 230058 13574 230614
rect 12954 194614 13574 230058
rect 16674 234334 17294 269778
rect 16674 233778 16706 234334
rect 17262 233778 17294 234334
rect 16208 219454 16528 219486
rect 16208 219218 16250 219454
rect 16486 219218 16528 219454
rect 16208 219134 16528 219218
rect 16208 218898 16250 219134
rect 16486 218898 16528 219134
rect 16208 218866 16528 218898
rect 12954 194058 12986 194614
rect 13542 194058 13574 194614
rect 12954 158614 13574 194058
rect 16674 198334 17294 233778
rect 16674 197778 16706 198334
rect 17262 197778 17294 198334
rect 16208 183454 16528 183486
rect 16208 183218 16250 183454
rect 16486 183218 16528 183454
rect 16208 183134 16528 183218
rect 16208 182898 16250 183134
rect 16486 182898 16528 183134
rect 16208 182866 16528 182898
rect 12954 158058 12986 158614
rect 13542 158058 13574 158614
rect 12954 122614 13574 158058
rect 16674 162334 17294 197778
rect 16674 161778 16706 162334
rect 17262 161778 17294 162334
rect 16208 147454 16528 147486
rect 16208 147218 16250 147454
rect 16486 147218 16528 147454
rect 16208 147134 16528 147218
rect 16208 146898 16250 147134
rect 16486 146898 16528 147134
rect 16208 146866 16528 146898
rect 12954 122058 12986 122614
rect 13542 122058 13574 122614
rect 12954 86614 13574 122058
rect 16674 126334 17294 161778
rect 16674 125778 16706 126334
rect 17262 125778 17294 126334
rect 16208 111454 16528 111486
rect 16208 111218 16250 111454
rect 16486 111218 16528 111454
rect 16208 111134 16528 111218
rect 16208 110898 16250 111134
rect 16486 110898 16528 111134
rect 16208 110866 16528 110898
rect 12954 86058 12986 86614
rect 13542 86058 13574 86614
rect 12954 50614 13574 86058
rect 16674 90334 17294 125778
rect 16674 89778 16706 90334
rect 17262 89778 17294 90334
rect 16208 75454 16528 75486
rect 16208 75218 16250 75454
rect 16486 75218 16528 75454
rect 16208 75134 16528 75218
rect 16208 74898 16250 75134
rect 16486 74898 16528 75134
rect 16208 74866 16528 74898
rect 12954 50058 12986 50614
rect 13542 50058 13574 50614
rect 12954 14614 13574 50058
rect 16674 54334 17294 89778
rect 16674 53778 16706 54334
rect 17262 53778 17294 54334
rect 16208 39454 16528 39486
rect 16208 39218 16250 39454
rect 16486 39218 16528 39454
rect 16208 39134 16528 39218
rect 16208 38898 16250 39134
rect 16486 38898 16528 39134
rect 16208 38866 16528 38898
rect 12954 14058 12986 14614
rect 13542 14058 13574 14614
rect 12954 -3226 13574 14058
rect 12954 -3782 12986 -3226
rect 13542 -3782 13574 -3226
rect 12954 -7654 13574 -3782
rect 16674 18334 17294 53778
rect 16674 17778 16706 18334
rect 17262 17778 17294 18334
rect 16674 -4186 17294 17778
rect 16674 -4742 16706 -4186
rect 17262 -4742 17294 -4186
rect 16674 -7654 17294 -4742
rect 20394 709638 21014 711590
rect 20394 709082 20426 709638
rect 20982 709082 21014 709638
rect 20394 670054 21014 709082
rect 20394 669498 20426 670054
rect 20982 669498 21014 670054
rect 20394 634054 21014 669498
rect 20394 633498 20426 634054
rect 20982 633498 21014 634054
rect 20394 598054 21014 633498
rect 20394 597498 20426 598054
rect 20982 597498 21014 598054
rect 20394 562054 21014 597498
rect 20394 561498 20426 562054
rect 20982 561498 21014 562054
rect 20394 526054 21014 561498
rect 20394 525498 20426 526054
rect 20982 525498 21014 526054
rect 20394 490054 21014 525498
rect 20394 489498 20426 490054
rect 20982 489498 21014 490054
rect 20394 454054 21014 489498
rect 20394 453498 20426 454054
rect 20982 453498 21014 454054
rect 20394 418054 21014 453498
rect 20394 417498 20426 418054
rect 20982 417498 21014 418054
rect 20394 382054 21014 417498
rect 20394 381498 20426 382054
rect 20982 381498 21014 382054
rect 20394 346054 21014 381498
rect 20394 345498 20426 346054
rect 20982 345498 21014 346054
rect 20394 310054 21014 345498
rect 20394 309498 20426 310054
rect 20982 309498 21014 310054
rect 20394 274054 21014 309498
rect 20394 273498 20426 274054
rect 20982 273498 21014 274054
rect 20394 238054 21014 273498
rect 20394 237498 20426 238054
rect 20982 237498 21014 238054
rect 20394 202054 21014 237498
rect 20394 201498 20426 202054
rect 20982 201498 21014 202054
rect 20394 166054 21014 201498
rect 20394 165498 20426 166054
rect 20982 165498 21014 166054
rect 20394 130054 21014 165498
rect 20394 129498 20426 130054
rect 20982 129498 21014 130054
rect 20394 94054 21014 129498
rect 20394 93498 20426 94054
rect 20982 93498 21014 94054
rect 20394 58054 21014 93498
rect 20394 57498 20426 58054
rect 20982 57498 21014 58054
rect 20394 22054 21014 57498
rect 20394 21498 20426 22054
rect 20982 21498 21014 22054
rect 20394 -5146 21014 21498
rect 20394 -5702 20426 -5146
rect 20982 -5702 21014 -5146
rect 20394 -7654 21014 -5702
rect 24114 710598 24734 711590
rect 24114 710042 24146 710598
rect 24702 710042 24734 710598
rect 24114 673774 24734 710042
rect 24114 673218 24146 673774
rect 24702 673218 24734 673774
rect 24114 637774 24734 673218
rect 24114 637218 24146 637774
rect 24702 637218 24734 637774
rect 24114 601774 24734 637218
rect 24114 601218 24146 601774
rect 24702 601218 24734 601774
rect 24114 565774 24734 601218
rect 24114 565218 24146 565774
rect 24702 565218 24734 565774
rect 24114 529774 24734 565218
rect 24114 529218 24146 529774
rect 24702 529218 24734 529774
rect 24114 493774 24734 529218
rect 24114 493218 24146 493774
rect 24702 493218 24734 493774
rect 24114 457774 24734 493218
rect 24114 457218 24146 457774
rect 24702 457218 24734 457774
rect 24114 421774 24734 457218
rect 24114 421218 24146 421774
rect 24702 421218 24734 421774
rect 24114 385774 24734 421218
rect 24114 385218 24146 385774
rect 24702 385218 24734 385774
rect 24114 349774 24734 385218
rect 24114 349218 24146 349774
rect 24702 349218 24734 349774
rect 24114 313774 24734 349218
rect 24114 313218 24146 313774
rect 24702 313218 24734 313774
rect 24114 277774 24734 313218
rect 24114 277218 24146 277774
rect 24702 277218 24734 277774
rect 24114 241774 24734 277218
rect 24114 241218 24146 241774
rect 24702 241218 24734 241774
rect 24114 205774 24734 241218
rect 24114 205218 24146 205774
rect 24702 205218 24734 205774
rect 24114 169774 24734 205218
rect 24114 169218 24146 169774
rect 24702 169218 24734 169774
rect 24114 133774 24734 169218
rect 24114 133218 24146 133774
rect 24702 133218 24734 133774
rect 24114 97774 24734 133218
rect 24114 97218 24146 97774
rect 24702 97218 24734 97774
rect 24114 61774 24734 97218
rect 24114 61218 24146 61774
rect 24702 61218 24734 61774
rect 24114 25774 24734 61218
rect 24114 25218 24146 25774
rect 24702 25218 24734 25774
rect 24114 -6106 24734 25218
rect 24114 -6662 24146 -6106
rect 24702 -6662 24734 -6106
rect 24114 -7654 24734 -6662
rect 27834 711558 28454 711590
rect 27834 711002 27866 711558
rect 28422 711002 28454 711558
rect 27834 677494 28454 711002
rect 27834 676938 27866 677494
rect 28422 676938 28454 677494
rect 27834 641494 28454 676938
rect 27834 640938 27866 641494
rect 28422 640938 28454 641494
rect 27834 605494 28454 640938
rect 27834 604938 27866 605494
rect 28422 604938 28454 605494
rect 27834 569494 28454 604938
rect 27834 568938 27866 569494
rect 28422 568938 28454 569494
rect 27834 533494 28454 568938
rect 27834 532938 27866 533494
rect 28422 532938 28454 533494
rect 27834 497494 28454 532938
rect 27834 496938 27866 497494
rect 28422 496938 28454 497494
rect 27834 461494 28454 496938
rect 27834 460938 27866 461494
rect 28422 460938 28454 461494
rect 27834 425494 28454 460938
rect 27834 424938 27866 425494
rect 28422 424938 28454 425494
rect 27834 389494 28454 424938
rect 27834 388938 27866 389494
rect 28422 388938 28454 389494
rect 27834 353494 28454 388938
rect 27834 352938 27866 353494
rect 28422 352938 28454 353494
rect 27834 317494 28454 352938
rect 37794 704838 38414 711590
rect 37794 704282 37826 704838
rect 38382 704282 38414 704838
rect 37794 687454 38414 704282
rect 37794 686898 37826 687454
rect 38382 686898 38414 687454
rect 37794 651454 38414 686898
rect 37794 650898 37826 651454
rect 38382 650898 38414 651454
rect 37794 615454 38414 650898
rect 37794 614898 37826 615454
rect 38382 614898 38414 615454
rect 37794 579454 38414 614898
rect 37794 578898 37826 579454
rect 38382 578898 38414 579454
rect 37794 543454 38414 578898
rect 37794 542898 37826 543454
rect 38382 542898 38414 543454
rect 37794 507454 38414 542898
rect 37794 506898 37826 507454
rect 38382 506898 38414 507454
rect 37794 471454 38414 506898
rect 37794 470898 37826 471454
rect 38382 470898 38414 471454
rect 37794 435454 38414 470898
rect 37794 434898 37826 435454
rect 38382 434898 38414 435454
rect 37794 399454 38414 434898
rect 37794 398898 37826 399454
rect 38382 398898 38414 399454
rect 37794 363454 38414 398898
rect 37794 362898 37826 363454
rect 38382 362898 38414 363454
rect 31568 331174 31888 331206
rect 31568 330938 31610 331174
rect 31846 330938 31888 331174
rect 31568 330854 31888 330938
rect 31568 330618 31610 330854
rect 31846 330618 31888 330854
rect 31568 330586 31888 330618
rect 27834 316938 27866 317494
rect 28422 316938 28454 317494
rect 27834 281494 28454 316938
rect 37794 327454 38414 362898
rect 37794 326898 37826 327454
rect 38382 326898 38414 327454
rect 31568 295174 31888 295206
rect 31568 294938 31610 295174
rect 31846 294938 31888 295174
rect 31568 294854 31888 294938
rect 31568 294618 31610 294854
rect 31846 294618 31888 294854
rect 31568 294586 31888 294618
rect 27834 280938 27866 281494
rect 28422 280938 28454 281494
rect 27834 245494 28454 280938
rect 37794 291454 38414 326898
rect 37794 290898 37826 291454
rect 38382 290898 38414 291454
rect 31568 259174 31888 259206
rect 31568 258938 31610 259174
rect 31846 258938 31888 259174
rect 31568 258854 31888 258938
rect 31568 258618 31610 258854
rect 31846 258618 31888 258854
rect 31568 258586 31888 258618
rect 27834 244938 27866 245494
rect 28422 244938 28454 245494
rect 27834 209494 28454 244938
rect 37794 255454 38414 290898
rect 37794 254898 37826 255454
rect 38382 254898 38414 255454
rect 31568 223174 31888 223206
rect 31568 222938 31610 223174
rect 31846 222938 31888 223174
rect 31568 222854 31888 222938
rect 31568 222618 31610 222854
rect 31846 222618 31888 222854
rect 31568 222586 31888 222618
rect 27834 208938 27866 209494
rect 28422 208938 28454 209494
rect 27834 173494 28454 208938
rect 37794 219454 38414 254898
rect 37794 218898 37826 219454
rect 38382 218898 38414 219454
rect 31568 187174 31888 187206
rect 31568 186938 31610 187174
rect 31846 186938 31888 187174
rect 31568 186854 31888 186938
rect 31568 186618 31610 186854
rect 31846 186618 31888 186854
rect 31568 186586 31888 186618
rect 27834 172938 27866 173494
rect 28422 172938 28454 173494
rect 27834 137494 28454 172938
rect 37794 183454 38414 218898
rect 37794 182898 37826 183454
rect 38382 182898 38414 183454
rect 31568 151174 31888 151206
rect 31568 150938 31610 151174
rect 31846 150938 31888 151174
rect 31568 150854 31888 150938
rect 31568 150618 31610 150854
rect 31846 150618 31888 150854
rect 31568 150586 31888 150618
rect 27834 136938 27866 137494
rect 28422 136938 28454 137494
rect 27834 101494 28454 136938
rect 37794 147454 38414 182898
rect 37794 146898 37826 147454
rect 38382 146898 38414 147454
rect 31568 115174 31888 115206
rect 31568 114938 31610 115174
rect 31846 114938 31888 115174
rect 31568 114854 31888 114938
rect 31568 114618 31610 114854
rect 31846 114618 31888 114854
rect 31568 114586 31888 114618
rect 27834 100938 27866 101494
rect 28422 100938 28454 101494
rect 27834 65494 28454 100938
rect 37794 111454 38414 146898
rect 37794 110898 37826 111454
rect 38382 110898 38414 111454
rect 31568 79174 31888 79206
rect 31568 78938 31610 79174
rect 31846 78938 31888 79174
rect 31568 78854 31888 78938
rect 31568 78618 31610 78854
rect 31846 78618 31888 78854
rect 31568 78586 31888 78618
rect 27834 64938 27866 65494
rect 28422 64938 28454 65494
rect 27834 29494 28454 64938
rect 37794 75454 38414 110898
rect 37794 74898 37826 75454
rect 38382 74898 38414 75454
rect 31568 43174 31888 43206
rect 31568 42938 31610 43174
rect 31846 42938 31888 43174
rect 31568 42854 31888 42938
rect 31568 42618 31610 42854
rect 31846 42618 31888 42854
rect 31568 42586 31888 42618
rect 27834 28938 27866 29494
rect 28422 28938 28454 29494
rect 27834 -7066 28454 28938
rect 37794 39454 38414 74898
rect 37794 38898 37826 39454
rect 38382 38898 38414 39454
rect 31568 7174 31888 7206
rect 31568 6938 31610 7174
rect 31846 6938 31888 7174
rect 31568 6854 31888 6938
rect 31568 6618 31610 6854
rect 31846 6618 31888 6854
rect 31568 6586 31888 6618
rect 27834 -7622 27866 -7066
rect 28422 -7622 28454 -7066
rect 27834 -7654 28454 -7622
rect 37794 3454 38414 38898
rect 37794 2898 37826 3454
rect 38382 2898 38414 3454
rect 37794 -346 38414 2898
rect 37794 -902 37826 -346
rect 38382 -902 38414 -346
rect 37794 -7654 38414 -902
rect 41514 705798 42134 711590
rect 41514 705242 41546 705798
rect 42102 705242 42134 705798
rect 41514 691174 42134 705242
rect 41514 690618 41546 691174
rect 42102 690618 42134 691174
rect 41514 655174 42134 690618
rect 41514 654618 41546 655174
rect 42102 654618 42134 655174
rect 41514 619174 42134 654618
rect 41514 618618 41546 619174
rect 42102 618618 42134 619174
rect 41514 583174 42134 618618
rect 41514 582618 41546 583174
rect 42102 582618 42134 583174
rect 41514 547174 42134 582618
rect 41514 546618 41546 547174
rect 42102 546618 42134 547174
rect 41514 511174 42134 546618
rect 41514 510618 41546 511174
rect 42102 510618 42134 511174
rect 41514 475174 42134 510618
rect 41514 474618 41546 475174
rect 42102 474618 42134 475174
rect 41514 439174 42134 474618
rect 41514 438618 41546 439174
rect 42102 438618 42134 439174
rect 41514 403174 42134 438618
rect 41514 402618 41546 403174
rect 42102 402618 42134 403174
rect 41514 367174 42134 402618
rect 41514 366618 41546 367174
rect 42102 366618 42134 367174
rect 41514 331174 42134 366618
rect 41514 330618 41546 331174
rect 42102 330618 42134 331174
rect 41514 295174 42134 330618
rect 41514 294618 41546 295174
rect 42102 294618 42134 295174
rect 41514 259174 42134 294618
rect 41514 258618 41546 259174
rect 42102 258618 42134 259174
rect 41514 223174 42134 258618
rect 41514 222618 41546 223174
rect 42102 222618 42134 223174
rect 41514 187174 42134 222618
rect 41514 186618 41546 187174
rect 42102 186618 42134 187174
rect 41514 151174 42134 186618
rect 41514 150618 41546 151174
rect 42102 150618 42134 151174
rect 41514 115174 42134 150618
rect 41514 114618 41546 115174
rect 42102 114618 42134 115174
rect 41514 79174 42134 114618
rect 41514 78618 41546 79174
rect 42102 78618 42134 79174
rect 41514 43174 42134 78618
rect 41514 42618 41546 43174
rect 42102 42618 42134 43174
rect 41514 7174 42134 42618
rect 41514 6618 41546 7174
rect 42102 6618 42134 7174
rect 41514 -1306 42134 6618
rect 41514 -1862 41546 -1306
rect 42102 -1862 42134 -1306
rect 41514 -7654 42134 -1862
rect 45234 706758 45854 711590
rect 45234 706202 45266 706758
rect 45822 706202 45854 706758
rect 45234 694894 45854 706202
rect 45234 694338 45266 694894
rect 45822 694338 45854 694894
rect 45234 658894 45854 694338
rect 45234 658338 45266 658894
rect 45822 658338 45854 658894
rect 45234 622894 45854 658338
rect 45234 622338 45266 622894
rect 45822 622338 45854 622894
rect 45234 586894 45854 622338
rect 45234 586338 45266 586894
rect 45822 586338 45854 586894
rect 45234 550894 45854 586338
rect 45234 550338 45266 550894
rect 45822 550338 45854 550894
rect 45234 514894 45854 550338
rect 45234 514338 45266 514894
rect 45822 514338 45854 514894
rect 45234 478894 45854 514338
rect 45234 478338 45266 478894
rect 45822 478338 45854 478894
rect 45234 442894 45854 478338
rect 45234 442338 45266 442894
rect 45822 442338 45854 442894
rect 45234 406894 45854 442338
rect 45234 406338 45266 406894
rect 45822 406338 45854 406894
rect 45234 370894 45854 406338
rect 45234 370338 45266 370894
rect 45822 370338 45854 370894
rect 45234 334894 45854 370338
rect 45234 334338 45266 334894
rect 45822 334338 45854 334894
rect 45234 298894 45854 334338
rect 48954 707718 49574 711590
rect 48954 707162 48986 707718
rect 49542 707162 49574 707718
rect 48954 698614 49574 707162
rect 48954 698058 48986 698614
rect 49542 698058 49574 698614
rect 48954 662614 49574 698058
rect 48954 662058 48986 662614
rect 49542 662058 49574 662614
rect 48954 626614 49574 662058
rect 48954 626058 48986 626614
rect 49542 626058 49574 626614
rect 48954 590614 49574 626058
rect 48954 590058 48986 590614
rect 49542 590058 49574 590614
rect 48954 554614 49574 590058
rect 48954 554058 48986 554614
rect 49542 554058 49574 554614
rect 48954 518614 49574 554058
rect 48954 518058 48986 518614
rect 49542 518058 49574 518614
rect 48954 482614 49574 518058
rect 48954 482058 48986 482614
rect 49542 482058 49574 482614
rect 48954 446614 49574 482058
rect 48954 446058 48986 446614
rect 49542 446058 49574 446614
rect 48954 410614 49574 446058
rect 48954 410058 48986 410614
rect 49542 410058 49574 410614
rect 48954 374614 49574 410058
rect 48954 374058 48986 374614
rect 49542 374058 49574 374614
rect 48954 338614 49574 374058
rect 48954 338058 48986 338614
rect 49542 338058 49574 338614
rect 46928 327454 47248 327486
rect 46928 327218 46970 327454
rect 47206 327218 47248 327454
rect 46928 327134 47248 327218
rect 46928 326898 46970 327134
rect 47206 326898 47248 327134
rect 46928 326866 47248 326898
rect 45234 298338 45266 298894
rect 45822 298338 45854 298894
rect 45234 262894 45854 298338
rect 48954 302614 49574 338058
rect 48954 302058 48986 302614
rect 49542 302058 49574 302614
rect 46928 291454 47248 291486
rect 46928 291218 46970 291454
rect 47206 291218 47248 291454
rect 46928 291134 47248 291218
rect 46928 290898 46970 291134
rect 47206 290898 47248 291134
rect 46928 290866 47248 290898
rect 45234 262338 45266 262894
rect 45822 262338 45854 262894
rect 45234 226894 45854 262338
rect 48954 266614 49574 302058
rect 48954 266058 48986 266614
rect 49542 266058 49574 266614
rect 46928 255454 47248 255486
rect 46928 255218 46970 255454
rect 47206 255218 47248 255454
rect 46928 255134 47248 255218
rect 46928 254898 46970 255134
rect 47206 254898 47248 255134
rect 46928 254866 47248 254898
rect 45234 226338 45266 226894
rect 45822 226338 45854 226894
rect 45234 190894 45854 226338
rect 48954 230614 49574 266058
rect 48954 230058 48986 230614
rect 49542 230058 49574 230614
rect 46928 219454 47248 219486
rect 46928 219218 46970 219454
rect 47206 219218 47248 219454
rect 46928 219134 47248 219218
rect 46928 218898 46970 219134
rect 47206 218898 47248 219134
rect 46928 218866 47248 218898
rect 45234 190338 45266 190894
rect 45822 190338 45854 190894
rect 45234 154894 45854 190338
rect 48954 194614 49574 230058
rect 48954 194058 48986 194614
rect 49542 194058 49574 194614
rect 46928 183454 47248 183486
rect 46928 183218 46970 183454
rect 47206 183218 47248 183454
rect 46928 183134 47248 183218
rect 46928 182898 46970 183134
rect 47206 182898 47248 183134
rect 46928 182866 47248 182898
rect 45234 154338 45266 154894
rect 45822 154338 45854 154894
rect 45234 118894 45854 154338
rect 48954 158614 49574 194058
rect 48954 158058 48986 158614
rect 49542 158058 49574 158614
rect 46928 147454 47248 147486
rect 46928 147218 46970 147454
rect 47206 147218 47248 147454
rect 46928 147134 47248 147218
rect 46928 146898 46970 147134
rect 47206 146898 47248 147134
rect 46928 146866 47248 146898
rect 45234 118338 45266 118894
rect 45822 118338 45854 118894
rect 45234 82894 45854 118338
rect 48954 122614 49574 158058
rect 48954 122058 48986 122614
rect 49542 122058 49574 122614
rect 46928 111454 47248 111486
rect 46928 111218 46970 111454
rect 47206 111218 47248 111454
rect 46928 111134 47248 111218
rect 46928 110898 46970 111134
rect 47206 110898 47248 111134
rect 46928 110866 47248 110898
rect 45234 82338 45266 82894
rect 45822 82338 45854 82894
rect 45234 46894 45854 82338
rect 48954 86614 49574 122058
rect 48954 86058 48986 86614
rect 49542 86058 49574 86614
rect 46928 75454 47248 75486
rect 46928 75218 46970 75454
rect 47206 75218 47248 75454
rect 46928 75134 47248 75218
rect 46928 74898 46970 75134
rect 47206 74898 47248 75134
rect 46928 74866 47248 74898
rect 45234 46338 45266 46894
rect 45822 46338 45854 46894
rect 45234 10894 45854 46338
rect 48954 50614 49574 86058
rect 48954 50058 48986 50614
rect 49542 50058 49574 50614
rect 46928 39454 47248 39486
rect 46928 39218 46970 39454
rect 47206 39218 47248 39454
rect 46928 39134 47248 39218
rect 46928 38898 46970 39134
rect 47206 38898 47248 39134
rect 46928 38866 47248 38898
rect 45234 10338 45266 10894
rect 45822 10338 45854 10894
rect 45234 -2266 45854 10338
rect 45234 -2822 45266 -2266
rect 45822 -2822 45854 -2266
rect 45234 -7654 45854 -2822
rect 48954 14614 49574 50058
rect 48954 14058 48986 14614
rect 49542 14058 49574 14614
rect 48954 -3226 49574 14058
rect 48954 -3782 48986 -3226
rect 49542 -3782 49574 -3226
rect 48954 -7654 49574 -3782
rect 52674 708678 53294 711590
rect 52674 708122 52706 708678
rect 53262 708122 53294 708678
rect 52674 666334 53294 708122
rect 52674 665778 52706 666334
rect 53262 665778 53294 666334
rect 52674 630334 53294 665778
rect 52674 629778 52706 630334
rect 53262 629778 53294 630334
rect 52674 594334 53294 629778
rect 52674 593778 52706 594334
rect 53262 593778 53294 594334
rect 52674 558334 53294 593778
rect 52674 557778 52706 558334
rect 53262 557778 53294 558334
rect 52674 522334 53294 557778
rect 52674 521778 52706 522334
rect 53262 521778 53294 522334
rect 52674 486334 53294 521778
rect 52674 485778 52706 486334
rect 53262 485778 53294 486334
rect 52674 450334 53294 485778
rect 52674 449778 52706 450334
rect 53262 449778 53294 450334
rect 52674 414334 53294 449778
rect 52674 413778 52706 414334
rect 53262 413778 53294 414334
rect 52674 378334 53294 413778
rect 52674 377778 52706 378334
rect 53262 377778 53294 378334
rect 52674 342334 53294 377778
rect 52674 341778 52706 342334
rect 53262 341778 53294 342334
rect 52674 306334 53294 341778
rect 52674 305778 52706 306334
rect 53262 305778 53294 306334
rect 52674 270334 53294 305778
rect 52674 269778 52706 270334
rect 53262 269778 53294 270334
rect 52674 234334 53294 269778
rect 52674 233778 52706 234334
rect 53262 233778 53294 234334
rect 52674 198334 53294 233778
rect 52674 197778 52706 198334
rect 53262 197778 53294 198334
rect 52674 162334 53294 197778
rect 52674 161778 52706 162334
rect 53262 161778 53294 162334
rect 52674 126334 53294 161778
rect 52674 125778 52706 126334
rect 53262 125778 53294 126334
rect 52674 90334 53294 125778
rect 52674 89778 52706 90334
rect 53262 89778 53294 90334
rect 52674 54334 53294 89778
rect 52674 53778 52706 54334
rect 53262 53778 53294 54334
rect 52674 18334 53294 53778
rect 52674 17778 52706 18334
rect 53262 17778 53294 18334
rect 52674 -4186 53294 17778
rect 52674 -4742 52706 -4186
rect 53262 -4742 53294 -4186
rect 52674 -7654 53294 -4742
rect 56394 709638 57014 711590
rect 56394 709082 56426 709638
rect 56982 709082 57014 709638
rect 56394 670054 57014 709082
rect 56394 669498 56426 670054
rect 56982 669498 57014 670054
rect 56394 634054 57014 669498
rect 56394 633498 56426 634054
rect 56982 633498 57014 634054
rect 56394 598054 57014 633498
rect 56394 597498 56426 598054
rect 56982 597498 57014 598054
rect 56394 562054 57014 597498
rect 56394 561498 56426 562054
rect 56982 561498 57014 562054
rect 56394 526054 57014 561498
rect 56394 525498 56426 526054
rect 56982 525498 57014 526054
rect 56394 490054 57014 525498
rect 56394 489498 56426 490054
rect 56982 489498 57014 490054
rect 56394 454054 57014 489498
rect 56394 453498 56426 454054
rect 56982 453498 57014 454054
rect 56394 418054 57014 453498
rect 56394 417498 56426 418054
rect 56982 417498 57014 418054
rect 56394 382054 57014 417498
rect 56394 381498 56426 382054
rect 56982 381498 57014 382054
rect 56394 346054 57014 381498
rect 56394 345498 56426 346054
rect 56982 345498 57014 346054
rect 56394 310054 57014 345498
rect 56394 309498 56426 310054
rect 56982 309498 57014 310054
rect 56394 274054 57014 309498
rect 56394 273498 56426 274054
rect 56982 273498 57014 274054
rect 56394 238054 57014 273498
rect 56394 237498 56426 238054
rect 56982 237498 57014 238054
rect 56394 202054 57014 237498
rect 56394 201498 56426 202054
rect 56982 201498 57014 202054
rect 56394 166054 57014 201498
rect 56394 165498 56426 166054
rect 56982 165498 57014 166054
rect 56394 130054 57014 165498
rect 56394 129498 56426 130054
rect 56982 129498 57014 130054
rect 56394 94054 57014 129498
rect 56394 93498 56426 94054
rect 56982 93498 57014 94054
rect 56394 58054 57014 93498
rect 56394 57498 56426 58054
rect 56982 57498 57014 58054
rect 56394 22054 57014 57498
rect 56394 21498 56426 22054
rect 56982 21498 57014 22054
rect 56394 -5146 57014 21498
rect 56394 -5702 56426 -5146
rect 56982 -5702 57014 -5146
rect 56394 -7654 57014 -5702
rect 60114 710598 60734 711590
rect 60114 710042 60146 710598
rect 60702 710042 60734 710598
rect 60114 673774 60734 710042
rect 60114 673218 60146 673774
rect 60702 673218 60734 673774
rect 60114 637774 60734 673218
rect 60114 637218 60146 637774
rect 60702 637218 60734 637774
rect 60114 601774 60734 637218
rect 60114 601218 60146 601774
rect 60702 601218 60734 601774
rect 60114 565774 60734 601218
rect 60114 565218 60146 565774
rect 60702 565218 60734 565774
rect 60114 529774 60734 565218
rect 60114 529218 60146 529774
rect 60702 529218 60734 529774
rect 60114 493774 60734 529218
rect 60114 493218 60146 493774
rect 60702 493218 60734 493774
rect 60114 457774 60734 493218
rect 60114 457218 60146 457774
rect 60702 457218 60734 457774
rect 60114 421774 60734 457218
rect 60114 421218 60146 421774
rect 60702 421218 60734 421774
rect 60114 385774 60734 421218
rect 60114 385218 60146 385774
rect 60702 385218 60734 385774
rect 60114 349774 60734 385218
rect 60114 349218 60146 349774
rect 60702 349218 60734 349774
rect 60114 313774 60734 349218
rect 63834 711558 64454 711590
rect 63834 711002 63866 711558
rect 64422 711002 64454 711558
rect 63834 677494 64454 711002
rect 63834 676938 63866 677494
rect 64422 676938 64454 677494
rect 63834 641494 64454 676938
rect 63834 640938 63866 641494
rect 64422 640938 64454 641494
rect 63834 605494 64454 640938
rect 63834 604938 63866 605494
rect 64422 604938 64454 605494
rect 63834 569494 64454 604938
rect 63834 568938 63866 569494
rect 64422 568938 64454 569494
rect 63834 533494 64454 568938
rect 63834 532938 63866 533494
rect 64422 532938 64454 533494
rect 63834 497494 64454 532938
rect 63834 496938 63866 497494
rect 64422 496938 64454 497494
rect 63834 461494 64454 496938
rect 63834 460938 63866 461494
rect 64422 460938 64454 461494
rect 63834 425494 64454 460938
rect 63834 424938 63866 425494
rect 64422 424938 64454 425494
rect 63834 389494 64454 424938
rect 63834 388938 63866 389494
rect 64422 388938 64454 389494
rect 63834 353494 64454 388938
rect 63834 352938 63866 353494
rect 64422 352938 64454 353494
rect 62288 331174 62608 331206
rect 62288 330938 62330 331174
rect 62566 330938 62608 331174
rect 62288 330854 62608 330938
rect 62288 330618 62330 330854
rect 62566 330618 62608 330854
rect 62288 330586 62608 330618
rect 60114 313218 60146 313774
rect 60702 313218 60734 313774
rect 60114 277774 60734 313218
rect 63834 317494 64454 352938
rect 63834 316938 63866 317494
rect 64422 316938 64454 317494
rect 62288 295174 62608 295206
rect 62288 294938 62330 295174
rect 62566 294938 62608 295174
rect 62288 294854 62608 294938
rect 62288 294618 62330 294854
rect 62566 294618 62608 294854
rect 62288 294586 62608 294618
rect 60114 277218 60146 277774
rect 60702 277218 60734 277774
rect 60114 241774 60734 277218
rect 63834 281494 64454 316938
rect 63834 280938 63866 281494
rect 64422 280938 64454 281494
rect 62288 259174 62608 259206
rect 62288 258938 62330 259174
rect 62566 258938 62608 259174
rect 62288 258854 62608 258938
rect 62288 258618 62330 258854
rect 62566 258618 62608 258854
rect 62288 258586 62608 258618
rect 60114 241218 60146 241774
rect 60702 241218 60734 241774
rect 60114 205774 60734 241218
rect 63834 245494 64454 280938
rect 63834 244938 63866 245494
rect 64422 244938 64454 245494
rect 62288 223174 62608 223206
rect 62288 222938 62330 223174
rect 62566 222938 62608 223174
rect 62288 222854 62608 222938
rect 62288 222618 62330 222854
rect 62566 222618 62608 222854
rect 62288 222586 62608 222618
rect 60114 205218 60146 205774
rect 60702 205218 60734 205774
rect 60114 169774 60734 205218
rect 63834 209494 64454 244938
rect 63834 208938 63866 209494
rect 64422 208938 64454 209494
rect 62288 187174 62608 187206
rect 62288 186938 62330 187174
rect 62566 186938 62608 187174
rect 62288 186854 62608 186938
rect 62288 186618 62330 186854
rect 62566 186618 62608 186854
rect 62288 186586 62608 186618
rect 60114 169218 60146 169774
rect 60702 169218 60734 169774
rect 60114 133774 60734 169218
rect 63834 173494 64454 208938
rect 63834 172938 63866 173494
rect 64422 172938 64454 173494
rect 62288 151174 62608 151206
rect 62288 150938 62330 151174
rect 62566 150938 62608 151174
rect 62288 150854 62608 150938
rect 62288 150618 62330 150854
rect 62566 150618 62608 150854
rect 62288 150586 62608 150618
rect 60114 133218 60146 133774
rect 60702 133218 60734 133774
rect 60114 97774 60734 133218
rect 63834 137494 64454 172938
rect 63834 136938 63866 137494
rect 64422 136938 64454 137494
rect 62288 115174 62608 115206
rect 62288 114938 62330 115174
rect 62566 114938 62608 115174
rect 62288 114854 62608 114938
rect 62288 114618 62330 114854
rect 62566 114618 62608 114854
rect 62288 114586 62608 114618
rect 60114 97218 60146 97774
rect 60702 97218 60734 97774
rect 60114 61774 60734 97218
rect 63834 101494 64454 136938
rect 63834 100938 63866 101494
rect 64422 100938 64454 101494
rect 62288 79174 62608 79206
rect 62288 78938 62330 79174
rect 62566 78938 62608 79174
rect 62288 78854 62608 78938
rect 62288 78618 62330 78854
rect 62566 78618 62608 78854
rect 62288 78586 62608 78618
rect 60114 61218 60146 61774
rect 60702 61218 60734 61774
rect 60114 25774 60734 61218
rect 63834 65494 64454 100938
rect 63834 64938 63866 65494
rect 64422 64938 64454 65494
rect 62288 43174 62608 43206
rect 62288 42938 62330 43174
rect 62566 42938 62608 43174
rect 62288 42854 62608 42938
rect 62288 42618 62330 42854
rect 62566 42618 62608 42854
rect 62288 42586 62608 42618
rect 60114 25218 60146 25774
rect 60702 25218 60734 25774
rect 60114 -6106 60734 25218
rect 63834 29494 64454 64938
rect 63834 28938 63866 29494
rect 64422 28938 64454 29494
rect 62288 7174 62608 7206
rect 62288 6938 62330 7174
rect 62566 6938 62608 7174
rect 62288 6854 62608 6938
rect 62288 6618 62330 6854
rect 62566 6618 62608 6854
rect 62288 6586 62608 6618
rect 60114 -6662 60146 -6106
rect 60702 -6662 60734 -6106
rect 60114 -7654 60734 -6662
rect 63834 -7066 64454 28938
rect 63834 -7622 63866 -7066
rect 64422 -7622 64454 -7066
rect 63834 -7654 64454 -7622
rect 73794 704838 74414 711590
rect 73794 704282 73826 704838
rect 74382 704282 74414 704838
rect 73794 687454 74414 704282
rect 73794 686898 73826 687454
rect 74382 686898 74414 687454
rect 73794 651454 74414 686898
rect 73794 650898 73826 651454
rect 74382 650898 74414 651454
rect 73794 615454 74414 650898
rect 73794 614898 73826 615454
rect 74382 614898 74414 615454
rect 73794 579454 74414 614898
rect 73794 578898 73826 579454
rect 74382 578898 74414 579454
rect 73794 543454 74414 578898
rect 73794 542898 73826 543454
rect 74382 542898 74414 543454
rect 73794 507454 74414 542898
rect 73794 506898 73826 507454
rect 74382 506898 74414 507454
rect 73794 471454 74414 506898
rect 73794 470898 73826 471454
rect 74382 470898 74414 471454
rect 73794 435454 74414 470898
rect 73794 434898 73826 435454
rect 74382 434898 74414 435454
rect 73794 399454 74414 434898
rect 73794 398898 73826 399454
rect 74382 398898 74414 399454
rect 73794 363454 74414 398898
rect 73794 362898 73826 363454
rect 74382 362898 74414 363454
rect 73794 327454 74414 362898
rect 77514 705798 78134 711590
rect 77514 705242 77546 705798
rect 78102 705242 78134 705798
rect 77514 691174 78134 705242
rect 77514 690618 77546 691174
rect 78102 690618 78134 691174
rect 77514 655174 78134 690618
rect 77514 654618 77546 655174
rect 78102 654618 78134 655174
rect 77514 619174 78134 654618
rect 77514 618618 77546 619174
rect 78102 618618 78134 619174
rect 77514 583174 78134 618618
rect 77514 582618 77546 583174
rect 78102 582618 78134 583174
rect 77514 547174 78134 582618
rect 77514 546618 77546 547174
rect 78102 546618 78134 547174
rect 77514 511174 78134 546618
rect 77514 510618 77546 511174
rect 78102 510618 78134 511174
rect 77514 475174 78134 510618
rect 77514 474618 77546 475174
rect 78102 474618 78134 475174
rect 77514 439174 78134 474618
rect 77514 438618 77546 439174
rect 78102 438618 78134 439174
rect 77514 403174 78134 438618
rect 77514 402618 77546 403174
rect 78102 402618 78134 403174
rect 77514 367174 78134 402618
rect 77514 366618 77546 367174
rect 78102 366618 78134 367174
rect 77514 354900 78134 366618
rect 81234 706758 81854 711590
rect 81234 706202 81266 706758
rect 81822 706202 81854 706758
rect 81234 694894 81854 706202
rect 81234 694338 81266 694894
rect 81822 694338 81854 694894
rect 81234 658894 81854 694338
rect 81234 658338 81266 658894
rect 81822 658338 81854 658894
rect 81234 622894 81854 658338
rect 81234 622338 81266 622894
rect 81822 622338 81854 622894
rect 81234 586894 81854 622338
rect 81234 586338 81266 586894
rect 81822 586338 81854 586894
rect 81234 550894 81854 586338
rect 81234 550338 81266 550894
rect 81822 550338 81854 550894
rect 81234 514894 81854 550338
rect 81234 514338 81266 514894
rect 81822 514338 81854 514894
rect 81234 478894 81854 514338
rect 81234 478338 81266 478894
rect 81822 478338 81854 478894
rect 81234 442894 81854 478338
rect 81234 442338 81266 442894
rect 81822 442338 81854 442894
rect 81234 406894 81854 442338
rect 81234 406338 81266 406894
rect 81822 406338 81854 406894
rect 81234 370894 81854 406338
rect 81234 370338 81266 370894
rect 81822 370338 81854 370894
rect 81234 334894 81854 370338
rect 81234 334338 81266 334894
rect 81822 334338 81854 334894
rect 73794 326898 73826 327454
rect 74382 326898 74414 327454
rect 73794 291454 74414 326898
rect 77648 327454 77968 327486
rect 77648 327218 77690 327454
rect 77926 327218 77968 327454
rect 77648 327134 77968 327218
rect 77648 326898 77690 327134
rect 77926 326898 77968 327134
rect 77648 326866 77968 326898
rect 81234 298894 81854 334338
rect 81234 298338 81266 298894
rect 81822 298338 81854 298894
rect 73794 290898 73826 291454
rect 74382 290898 74414 291454
rect 73794 255454 74414 290898
rect 77648 291454 77968 291486
rect 77648 291218 77690 291454
rect 77926 291218 77968 291454
rect 77648 291134 77968 291218
rect 77648 290898 77690 291134
rect 77926 290898 77968 291134
rect 77648 290866 77968 290898
rect 81234 262894 81854 298338
rect 81234 262338 81266 262894
rect 81822 262338 81854 262894
rect 73794 254898 73826 255454
rect 74382 254898 74414 255454
rect 73794 219454 74414 254898
rect 77648 255454 77968 255486
rect 77648 255218 77690 255454
rect 77926 255218 77968 255454
rect 77648 255134 77968 255218
rect 77648 254898 77690 255134
rect 77926 254898 77968 255134
rect 77648 254866 77968 254898
rect 81234 226894 81854 262338
rect 81234 226338 81266 226894
rect 81822 226338 81854 226894
rect 73794 218898 73826 219454
rect 74382 218898 74414 219454
rect 73794 183454 74414 218898
rect 77648 219454 77968 219486
rect 77648 219218 77690 219454
rect 77926 219218 77968 219454
rect 77648 219134 77968 219218
rect 77648 218898 77690 219134
rect 77926 218898 77968 219134
rect 77648 218866 77968 218898
rect 81234 190894 81854 226338
rect 81234 190338 81266 190894
rect 81822 190338 81854 190894
rect 73794 182898 73826 183454
rect 74382 182898 74414 183454
rect 73794 147454 74414 182898
rect 77648 183454 77968 183486
rect 77648 183218 77690 183454
rect 77926 183218 77968 183454
rect 77648 183134 77968 183218
rect 77648 182898 77690 183134
rect 77926 182898 77968 183134
rect 77648 182866 77968 182898
rect 81234 154894 81854 190338
rect 81234 154338 81266 154894
rect 81822 154338 81854 154894
rect 73794 146898 73826 147454
rect 74382 146898 74414 147454
rect 73794 111454 74414 146898
rect 77648 147454 77968 147486
rect 77648 147218 77690 147454
rect 77926 147218 77968 147454
rect 77648 147134 77968 147218
rect 77648 146898 77690 147134
rect 77926 146898 77968 147134
rect 77648 146866 77968 146898
rect 81234 118894 81854 154338
rect 81234 118338 81266 118894
rect 81822 118338 81854 118894
rect 73794 110898 73826 111454
rect 74382 110898 74414 111454
rect 73794 75454 74414 110898
rect 77648 111454 77968 111486
rect 77648 111218 77690 111454
rect 77926 111218 77968 111454
rect 77648 111134 77968 111218
rect 77648 110898 77690 111134
rect 77926 110898 77968 111134
rect 77648 110866 77968 110898
rect 81234 82894 81854 118338
rect 81234 82338 81266 82894
rect 81822 82338 81854 82894
rect 73794 74898 73826 75454
rect 74382 74898 74414 75454
rect 73794 39454 74414 74898
rect 77648 75454 77968 75486
rect 77648 75218 77690 75454
rect 77926 75218 77968 75454
rect 77648 75134 77968 75218
rect 77648 74898 77690 75134
rect 77926 74898 77968 75134
rect 77648 74866 77968 74898
rect 81234 46894 81854 82338
rect 81234 46338 81266 46894
rect 81822 46338 81854 46894
rect 73794 38898 73826 39454
rect 74382 38898 74414 39454
rect 73794 3454 74414 38898
rect 77648 39454 77968 39486
rect 77648 39218 77690 39454
rect 77926 39218 77968 39454
rect 77648 39134 77968 39218
rect 77648 38898 77690 39134
rect 77926 38898 77968 39134
rect 77648 38866 77968 38898
rect 73794 2898 73826 3454
rect 74382 2898 74414 3454
rect 73794 -346 74414 2898
rect 73794 -902 73826 -346
rect 74382 -902 74414 -346
rect 73794 -7654 74414 -902
rect 81234 10894 81854 46338
rect 81234 10338 81266 10894
rect 81822 10338 81854 10894
rect 81234 -2266 81854 10338
rect 81234 -2822 81266 -2266
rect 81822 -2822 81854 -2266
rect 81234 -7654 81854 -2822
rect 84954 707718 85574 711590
rect 84954 707162 84986 707718
rect 85542 707162 85574 707718
rect 84954 698614 85574 707162
rect 84954 698058 84986 698614
rect 85542 698058 85574 698614
rect 84954 662614 85574 698058
rect 84954 662058 84986 662614
rect 85542 662058 85574 662614
rect 84954 626614 85574 662058
rect 84954 626058 84986 626614
rect 85542 626058 85574 626614
rect 84954 590614 85574 626058
rect 84954 590058 84986 590614
rect 85542 590058 85574 590614
rect 84954 554614 85574 590058
rect 84954 554058 84986 554614
rect 85542 554058 85574 554614
rect 84954 518614 85574 554058
rect 84954 518058 84986 518614
rect 85542 518058 85574 518614
rect 84954 482614 85574 518058
rect 84954 482058 84986 482614
rect 85542 482058 85574 482614
rect 84954 446614 85574 482058
rect 84954 446058 84986 446614
rect 85542 446058 85574 446614
rect 84954 410614 85574 446058
rect 84954 410058 84986 410614
rect 85542 410058 85574 410614
rect 84954 374614 85574 410058
rect 84954 374058 84986 374614
rect 85542 374058 85574 374614
rect 84954 338614 85574 374058
rect 84954 338058 84986 338614
rect 85542 338058 85574 338614
rect 84954 302614 85574 338058
rect 84954 302058 84986 302614
rect 85542 302058 85574 302614
rect 84954 266614 85574 302058
rect 84954 266058 84986 266614
rect 85542 266058 85574 266614
rect 84954 230614 85574 266058
rect 84954 230058 84986 230614
rect 85542 230058 85574 230614
rect 84954 194614 85574 230058
rect 84954 194058 84986 194614
rect 85542 194058 85574 194614
rect 84954 158614 85574 194058
rect 84954 158058 84986 158614
rect 85542 158058 85574 158614
rect 84954 122614 85574 158058
rect 84954 122058 84986 122614
rect 85542 122058 85574 122614
rect 84954 86614 85574 122058
rect 84954 86058 84986 86614
rect 85542 86058 85574 86614
rect 84954 50614 85574 86058
rect 84954 50058 84986 50614
rect 85542 50058 85574 50614
rect 84954 14614 85574 50058
rect 84954 14058 84986 14614
rect 85542 14058 85574 14614
rect 84954 -3226 85574 14058
rect 84954 -3782 84986 -3226
rect 85542 -3782 85574 -3226
rect 84954 -7654 85574 -3782
rect 88674 708678 89294 711590
rect 88674 708122 88706 708678
rect 89262 708122 89294 708678
rect 88674 666334 89294 708122
rect 88674 665778 88706 666334
rect 89262 665778 89294 666334
rect 88674 630334 89294 665778
rect 88674 629778 88706 630334
rect 89262 629778 89294 630334
rect 88674 594334 89294 629778
rect 88674 593778 88706 594334
rect 89262 593778 89294 594334
rect 88674 558334 89294 593778
rect 88674 557778 88706 558334
rect 89262 557778 89294 558334
rect 88674 522334 89294 557778
rect 88674 521778 88706 522334
rect 89262 521778 89294 522334
rect 88674 486334 89294 521778
rect 88674 485778 88706 486334
rect 89262 485778 89294 486334
rect 88674 450334 89294 485778
rect 88674 449778 88706 450334
rect 89262 449778 89294 450334
rect 88674 414334 89294 449778
rect 88674 413778 88706 414334
rect 89262 413778 89294 414334
rect 88674 378334 89294 413778
rect 88674 377778 88706 378334
rect 89262 377778 89294 378334
rect 88674 342334 89294 377778
rect 92394 709638 93014 711590
rect 92394 709082 92426 709638
rect 92982 709082 93014 709638
rect 92394 670054 93014 709082
rect 92394 669498 92426 670054
rect 92982 669498 93014 670054
rect 92394 634054 93014 669498
rect 92394 633498 92426 634054
rect 92982 633498 93014 634054
rect 92394 598054 93014 633498
rect 92394 597498 92426 598054
rect 92982 597498 93014 598054
rect 92394 562054 93014 597498
rect 92394 561498 92426 562054
rect 92982 561498 93014 562054
rect 92394 526054 93014 561498
rect 92394 525498 92426 526054
rect 92982 525498 93014 526054
rect 92394 490054 93014 525498
rect 92394 489498 92426 490054
rect 92982 489498 93014 490054
rect 92394 454054 93014 489498
rect 92394 453498 92426 454054
rect 92982 453498 93014 454054
rect 92394 418054 93014 453498
rect 92394 417498 92426 418054
rect 92982 417498 93014 418054
rect 92394 382054 93014 417498
rect 92394 381498 92426 382054
rect 92982 381498 93014 382054
rect 92394 354900 93014 381498
rect 96114 710598 96734 711590
rect 96114 710042 96146 710598
rect 96702 710042 96734 710598
rect 96114 673774 96734 710042
rect 96114 673218 96146 673774
rect 96702 673218 96734 673774
rect 96114 637774 96734 673218
rect 96114 637218 96146 637774
rect 96702 637218 96734 637774
rect 96114 601774 96734 637218
rect 96114 601218 96146 601774
rect 96702 601218 96734 601774
rect 96114 565774 96734 601218
rect 96114 565218 96146 565774
rect 96702 565218 96734 565774
rect 96114 529774 96734 565218
rect 96114 529218 96146 529774
rect 96702 529218 96734 529774
rect 96114 493774 96734 529218
rect 96114 493218 96146 493774
rect 96702 493218 96734 493774
rect 96114 457774 96734 493218
rect 96114 457218 96146 457774
rect 96702 457218 96734 457774
rect 96114 421774 96734 457218
rect 96114 421218 96146 421774
rect 96702 421218 96734 421774
rect 96114 385774 96734 421218
rect 96114 385218 96146 385774
rect 96702 385218 96734 385774
rect 88674 341778 88706 342334
rect 89262 341778 89294 342334
rect 88674 306334 89294 341778
rect 96114 349774 96734 385218
rect 96114 349218 96146 349774
rect 96702 349218 96734 349774
rect 93008 331174 93328 331206
rect 93008 330938 93050 331174
rect 93286 330938 93328 331174
rect 93008 330854 93328 330938
rect 93008 330618 93050 330854
rect 93286 330618 93328 330854
rect 93008 330586 93328 330618
rect 88674 305778 88706 306334
rect 89262 305778 89294 306334
rect 88674 270334 89294 305778
rect 96114 313774 96734 349218
rect 96114 313218 96146 313774
rect 96702 313218 96734 313774
rect 93008 295174 93328 295206
rect 93008 294938 93050 295174
rect 93286 294938 93328 295174
rect 93008 294854 93328 294938
rect 93008 294618 93050 294854
rect 93286 294618 93328 294854
rect 93008 294586 93328 294618
rect 88674 269778 88706 270334
rect 89262 269778 89294 270334
rect 88674 234334 89294 269778
rect 96114 277774 96734 313218
rect 96114 277218 96146 277774
rect 96702 277218 96734 277774
rect 93008 259174 93328 259206
rect 93008 258938 93050 259174
rect 93286 258938 93328 259174
rect 93008 258854 93328 258938
rect 93008 258618 93050 258854
rect 93286 258618 93328 258854
rect 93008 258586 93328 258618
rect 88674 233778 88706 234334
rect 89262 233778 89294 234334
rect 88674 198334 89294 233778
rect 96114 241774 96734 277218
rect 96114 241218 96146 241774
rect 96702 241218 96734 241774
rect 93008 223174 93328 223206
rect 93008 222938 93050 223174
rect 93286 222938 93328 223174
rect 93008 222854 93328 222938
rect 93008 222618 93050 222854
rect 93286 222618 93328 222854
rect 93008 222586 93328 222618
rect 88674 197778 88706 198334
rect 89262 197778 89294 198334
rect 88674 162334 89294 197778
rect 96114 205774 96734 241218
rect 96114 205218 96146 205774
rect 96702 205218 96734 205774
rect 93008 187174 93328 187206
rect 93008 186938 93050 187174
rect 93286 186938 93328 187174
rect 93008 186854 93328 186938
rect 93008 186618 93050 186854
rect 93286 186618 93328 186854
rect 93008 186586 93328 186618
rect 88674 161778 88706 162334
rect 89262 161778 89294 162334
rect 88674 126334 89294 161778
rect 96114 169774 96734 205218
rect 96114 169218 96146 169774
rect 96702 169218 96734 169774
rect 93008 151174 93328 151206
rect 93008 150938 93050 151174
rect 93286 150938 93328 151174
rect 93008 150854 93328 150938
rect 93008 150618 93050 150854
rect 93286 150618 93328 150854
rect 93008 150586 93328 150618
rect 88674 125778 88706 126334
rect 89262 125778 89294 126334
rect 88674 90334 89294 125778
rect 96114 133774 96734 169218
rect 96114 133218 96146 133774
rect 96702 133218 96734 133774
rect 93008 115174 93328 115206
rect 93008 114938 93050 115174
rect 93286 114938 93328 115174
rect 93008 114854 93328 114938
rect 93008 114618 93050 114854
rect 93286 114618 93328 114854
rect 93008 114586 93328 114618
rect 88674 89778 88706 90334
rect 89262 89778 89294 90334
rect 88674 54334 89294 89778
rect 96114 97774 96734 133218
rect 96114 97218 96146 97774
rect 96702 97218 96734 97774
rect 93008 79174 93328 79206
rect 93008 78938 93050 79174
rect 93286 78938 93328 79174
rect 93008 78854 93328 78938
rect 93008 78618 93050 78854
rect 93286 78618 93328 78854
rect 93008 78586 93328 78618
rect 88674 53778 88706 54334
rect 89262 53778 89294 54334
rect 88674 18334 89294 53778
rect 96114 61774 96734 97218
rect 96114 61218 96146 61774
rect 96702 61218 96734 61774
rect 93008 43174 93328 43206
rect 93008 42938 93050 43174
rect 93286 42938 93328 43174
rect 93008 42854 93328 42938
rect 93008 42618 93050 42854
rect 93286 42618 93328 42854
rect 93008 42586 93328 42618
rect 88674 17778 88706 18334
rect 89262 17778 89294 18334
rect 88674 -4186 89294 17778
rect 96114 25774 96734 61218
rect 96114 25218 96146 25774
rect 96702 25218 96734 25774
rect 93008 7174 93328 7206
rect 93008 6938 93050 7174
rect 93286 6938 93328 7174
rect 93008 6854 93328 6938
rect 93008 6618 93050 6854
rect 93286 6618 93328 6854
rect 93008 6586 93328 6618
rect 88674 -4742 88706 -4186
rect 89262 -4742 89294 -4186
rect 88674 -7654 89294 -4742
rect 96114 -6106 96734 25218
rect 96114 -6662 96146 -6106
rect 96702 -6662 96734 -6106
rect 96114 -7654 96734 -6662
rect 99834 711558 100454 711590
rect 99834 711002 99866 711558
rect 100422 711002 100454 711558
rect 99834 677494 100454 711002
rect 99834 676938 99866 677494
rect 100422 676938 100454 677494
rect 99834 641494 100454 676938
rect 99834 640938 99866 641494
rect 100422 640938 100454 641494
rect 99834 605494 100454 640938
rect 99834 604938 99866 605494
rect 100422 604938 100454 605494
rect 99834 569494 100454 604938
rect 99834 568938 99866 569494
rect 100422 568938 100454 569494
rect 99834 533494 100454 568938
rect 99834 532938 99866 533494
rect 100422 532938 100454 533494
rect 99834 497494 100454 532938
rect 99834 496938 99866 497494
rect 100422 496938 100454 497494
rect 99834 461494 100454 496938
rect 99834 460938 99866 461494
rect 100422 460938 100454 461494
rect 99834 425494 100454 460938
rect 99834 424938 99866 425494
rect 100422 424938 100454 425494
rect 99834 389494 100454 424938
rect 99834 388938 99866 389494
rect 100422 388938 100454 389494
rect 99834 353494 100454 388938
rect 99834 352938 99866 353494
rect 100422 352938 100454 353494
rect 99834 317494 100454 352938
rect 109794 704838 110414 711590
rect 109794 704282 109826 704838
rect 110382 704282 110414 704838
rect 109794 687454 110414 704282
rect 109794 686898 109826 687454
rect 110382 686898 110414 687454
rect 109794 651454 110414 686898
rect 109794 650898 109826 651454
rect 110382 650898 110414 651454
rect 109794 615454 110414 650898
rect 109794 614898 109826 615454
rect 110382 614898 110414 615454
rect 109794 579454 110414 614898
rect 109794 578898 109826 579454
rect 110382 578898 110414 579454
rect 109794 543454 110414 578898
rect 109794 542898 109826 543454
rect 110382 542898 110414 543454
rect 109794 507454 110414 542898
rect 109794 506898 109826 507454
rect 110382 506898 110414 507454
rect 109794 471454 110414 506898
rect 109794 470898 109826 471454
rect 110382 470898 110414 471454
rect 109794 435454 110414 470898
rect 109794 434898 109826 435454
rect 110382 434898 110414 435454
rect 109794 399454 110414 434898
rect 109794 398898 109826 399454
rect 110382 398898 110414 399454
rect 109794 363454 110414 398898
rect 109794 362898 109826 363454
rect 110382 362898 110414 363454
rect 108368 327454 108688 327486
rect 108368 327218 108410 327454
rect 108646 327218 108688 327454
rect 108368 327134 108688 327218
rect 108368 326898 108410 327134
rect 108646 326898 108688 327134
rect 108368 326866 108688 326898
rect 109794 327454 110414 362898
rect 109794 326898 109826 327454
rect 110382 326898 110414 327454
rect 99834 316938 99866 317494
rect 100422 316938 100454 317494
rect 99834 281494 100454 316938
rect 108368 291454 108688 291486
rect 108368 291218 108410 291454
rect 108646 291218 108688 291454
rect 108368 291134 108688 291218
rect 108368 290898 108410 291134
rect 108646 290898 108688 291134
rect 108368 290866 108688 290898
rect 109794 291454 110414 326898
rect 109794 290898 109826 291454
rect 110382 290898 110414 291454
rect 99834 280938 99866 281494
rect 100422 280938 100454 281494
rect 99834 245494 100454 280938
rect 108368 255454 108688 255486
rect 108368 255218 108410 255454
rect 108646 255218 108688 255454
rect 108368 255134 108688 255218
rect 108368 254898 108410 255134
rect 108646 254898 108688 255134
rect 108368 254866 108688 254898
rect 109794 255454 110414 290898
rect 109794 254898 109826 255454
rect 110382 254898 110414 255454
rect 99834 244938 99866 245494
rect 100422 244938 100454 245494
rect 99834 209494 100454 244938
rect 108368 219454 108688 219486
rect 108368 219218 108410 219454
rect 108646 219218 108688 219454
rect 108368 219134 108688 219218
rect 108368 218898 108410 219134
rect 108646 218898 108688 219134
rect 108368 218866 108688 218898
rect 109794 219454 110414 254898
rect 109794 218898 109826 219454
rect 110382 218898 110414 219454
rect 99834 208938 99866 209494
rect 100422 208938 100454 209494
rect 99834 173494 100454 208938
rect 108368 183454 108688 183486
rect 108368 183218 108410 183454
rect 108646 183218 108688 183454
rect 108368 183134 108688 183218
rect 108368 182898 108410 183134
rect 108646 182898 108688 183134
rect 108368 182866 108688 182898
rect 109794 183454 110414 218898
rect 109794 182898 109826 183454
rect 110382 182898 110414 183454
rect 99834 172938 99866 173494
rect 100422 172938 100454 173494
rect 99834 137494 100454 172938
rect 108368 147454 108688 147486
rect 108368 147218 108410 147454
rect 108646 147218 108688 147454
rect 108368 147134 108688 147218
rect 108368 146898 108410 147134
rect 108646 146898 108688 147134
rect 108368 146866 108688 146898
rect 109794 147454 110414 182898
rect 109794 146898 109826 147454
rect 110382 146898 110414 147454
rect 99834 136938 99866 137494
rect 100422 136938 100454 137494
rect 99834 101494 100454 136938
rect 108368 111454 108688 111486
rect 108368 111218 108410 111454
rect 108646 111218 108688 111454
rect 108368 111134 108688 111218
rect 108368 110898 108410 111134
rect 108646 110898 108688 111134
rect 108368 110866 108688 110898
rect 109794 111454 110414 146898
rect 109794 110898 109826 111454
rect 110382 110898 110414 111454
rect 99834 100938 99866 101494
rect 100422 100938 100454 101494
rect 99834 65494 100454 100938
rect 108368 75454 108688 75486
rect 108368 75218 108410 75454
rect 108646 75218 108688 75454
rect 108368 75134 108688 75218
rect 108368 74898 108410 75134
rect 108646 74898 108688 75134
rect 108368 74866 108688 74898
rect 109794 75454 110414 110898
rect 109794 74898 109826 75454
rect 110382 74898 110414 75454
rect 99834 64938 99866 65494
rect 100422 64938 100454 65494
rect 99834 29494 100454 64938
rect 108368 39454 108688 39486
rect 108368 39218 108410 39454
rect 108646 39218 108688 39454
rect 108368 39134 108688 39218
rect 108368 38898 108410 39134
rect 108646 38898 108688 39134
rect 108368 38866 108688 38898
rect 109794 39454 110414 74898
rect 109794 38898 109826 39454
rect 110382 38898 110414 39454
rect 99834 28938 99866 29494
rect 100422 28938 100454 29494
rect 99834 -7066 100454 28938
rect 99834 -7622 99866 -7066
rect 100422 -7622 100454 -7066
rect 99834 -7654 100454 -7622
rect 109794 3454 110414 38898
rect 109794 2898 109826 3454
rect 110382 2898 110414 3454
rect 109794 -346 110414 2898
rect 109794 -902 109826 -346
rect 110382 -902 110414 -346
rect 109794 -7654 110414 -902
rect 113514 705798 114134 711590
rect 113514 705242 113546 705798
rect 114102 705242 114134 705798
rect 113514 691174 114134 705242
rect 113514 690618 113546 691174
rect 114102 690618 114134 691174
rect 113514 655174 114134 690618
rect 113514 654618 113546 655174
rect 114102 654618 114134 655174
rect 113514 619174 114134 654618
rect 113514 618618 113546 619174
rect 114102 618618 114134 619174
rect 113514 583174 114134 618618
rect 113514 582618 113546 583174
rect 114102 582618 114134 583174
rect 113514 547174 114134 582618
rect 113514 546618 113546 547174
rect 114102 546618 114134 547174
rect 113514 511174 114134 546618
rect 113514 510618 113546 511174
rect 114102 510618 114134 511174
rect 113514 475174 114134 510618
rect 113514 474618 113546 475174
rect 114102 474618 114134 475174
rect 113514 439174 114134 474618
rect 113514 438618 113546 439174
rect 114102 438618 114134 439174
rect 113514 403174 114134 438618
rect 113514 402618 113546 403174
rect 114102 402618 114134 403174
rect 113514 367174 114134 402618
rect 113514 366618 113546 367174
rect 114102 366618 114134 367174
rect 113514 331174 114134 366618
rect 113514 330618 113546 331174
rect 114102 330618 114134 331174
rect 113514 295174 114134 330618
rect 113514 294618 113546 295174
rect 114102 294618 114134 295174
rect 113514 259174 114134 294618
rect 113514 258618 113546 259174
rect 114102 258618 114134 259174
rect 113514 223174 114134 258618
rect 113514 222618 113546 223174
rect 114102 222618 114134 223174
rect 113514 187174 114134 222618
rect 113514 186618 113546 187174
rect 114102 186618 114134 187174
rect 113514 151174 114134 186618
rect 113514 150618 113546 151174
rect 114102 150618 114134 151174
rect 113514 115174 114134 150618
rect 113514 114618 113546 115174
rect 114102 114618 114134 115174
rect 113514 79174 114134 114618
rect 113514 78618 113546 79174
rect 114102 78618 114134 79174
rect 113514 43174 114134 78618
rect 113514 42618 113546 43174
rect 114102 42618 114134 43174
rect 113514 7174 114134 42618
rect 113514 6618 113546 7174
rect 114102 6618 114134 7174
rect 113514 -1306 114134 6618
rect 113514 -1862 113546 -1306
rect 114102 -1862 114134 -1306
rect 113514 -7654 114134 -1862
rect 117234 706758 117854 711590
rect 117234 706202 117266 706758
rect 117822 706202 117854 706758
rect 117234 694894 117854 706202
rect 117234 694338 117266 694894
rect 117822 694338 117854 694894
rect 117234 658894 117854 694338
rect 117234 658338 117266 658894
rect 117822 658338 117854 658894
rect 117234 622894 117854 658338
rect 117234 622338 117266 622894
rect 117822 622338 117854 622894
rect 117234 586894 117854 622338
rect 117234 586338 117266 586894
rect 117822 586338 117854 586894
rect 117234 550894 117854 586338
rect 117234 550338 117266 550894
rect 117822 550338 117854 550894
rect 117234 514894 117854 550338
rect 117234 514338 117266 514894
rect 117822 514338 117854 514894
rect 117234 478894 117854 514338
rect 117234 478338 117266 478894
rect 117822 478338 117854 478894
rect 117234 442894 117854 478338
rect 117234 442338 117266 442894
rect 117822 442338 117854 442894
rect 117234 406894 117854 442338
rect 117234 406338 117266 406894
rect 117822 406338 117854 406894
rect 117234 370894 117854 406338
rect 117234 370338 117266 370894
rect 117822 370338 117854 370894
rect 117234 334894 117854 370338
rect 117234 334338 117266 334894
rect 117822 334338 117854 334894
rect 117234 298894 117854 334338
rect 117234 298338 117266 298894
rect 117822 298338 117854 298894
rect 117234 262894 117854 298338
rect 117234 262338 117266 262894
rect 117822 262338 117854 262894
rect 117234 226894 117854 262338
rect 117234 226338 117266 226894
rect 117822 226338 117854 226894
rect 117234 190894 117854 226338
rect 117234 190338 117266 190894
rect 117822 190338 117854 190894
rect 117234 154894 117854 190338
rect 117234 154338 117266 154894
rect 117822 154338 117854 154894
rect 117234 118894 117854 154338
rect 117234 118338 117266 118894
rect 117822 118338 117854 118894
rect 117234 82894 117854 118338
rect 117234 82338 117266 82894
rect 117822 82338 117854 82894
rect 117234 46894 117854 82338
rect 117234 46338 117266 46894
rect 117822 46338 117854 46894
rect 117234 10894 117854 46338
rect 117234 10338 117266 10894
rect 117822 10338 117854 10894
rect 117234 -2266 117854 10338
rect 117234 -2822 117266 -2266
rect 117822 -2822 117854 -2266
rect 117234 -7654 117854 -2822
rect 120954 707718 121574 711590
rect 120954 707162 120986 707718
rect 121542 707162 121574 707718
rect 120954 698614 121574 707162
rect 120954 698058 120986 698614
rect 121542 698058 121574 698614
rect 120954 662614 121574 698058
rect 120954 662058 120986 662614
rect 121542 662058 121574 662614
rect 120954 626614 121574 662058
rect 120954 626058 120986 626614
rect 121542 626058 121574 626614
rect 120954 590614 121574 626058
rect 120954 590058 120986 590614
rect 121542 590058 121574 590614
rect 120954 554614 121574 590058
rect 120954 554058 120986 554614
rect 121542 554058 121574 554614
rect 120954 518614 121574 554058
rect 120954 518058 120986 518614
rect 121542 518058 121574 518614
rect 120954 482614 121574 518058
rect 120954 482058 120986 482614
rect 121542 482058 121574 482614
rect 120954 446614 121574 482058
rect 120954 446058 120986 446614
rect 121542 446058 121574 446614
rect 120954 410614 121574 446058
rect 120954 410058 120986 410614
rect 121542 410058 121574 410614
rect 120954 374614 121574 410058
rect 120954 374058 120986 374614
rect 121542 374058 121574 374614
rect 120954 338614 121574 374058
rect 120954 338058 120986 338614
rect 121542 338058 121574 338614
rect 120954 302614 121574 338058
rect 124674 708678 125294 711590
rect 124674 708122 124706 708678
rect 125262 708122 125294 708678
rect 124674 666334 125294 708122
rect 124674 665778 124706 666334
rect 125262 665778 125294 666334
rect 124674 630334 125294 665778
rect 124674 629778 124706 630334
rect 125262 629778 125294 630334
rect 124674 594334 125294 629778
rect 124674 593778 124706 594334
rect 125262 593778 125294 594334
rect 124674 558334 125294 593778
rect 124674 557778 124706 558334
rect 125262 557778 125294 558334
rect 124674 522334 125294 557778
rect 124674 521778 124706 522334
rect 125262 521778 125294 522334
rect 124674 486334 125294 521778
rect 124674 485778 124706 486334
rect 125262 485778 125294 486334
rect 124674 450334 125294 485778
rect 124674 449778 124706 450334
rect 125262 449778 125294 450334
rect 124674 414334 125294 449778
rect 124674 413778 124706 414334
rect 125262 413778 125294 414334
rect 124674 378334 125294 413778
rect 124674 377778 124706 378334
rect 125262 377778 125294 378334
rect 124674 342334 125294 377778
rect 124674 341778 124706 342334
rect 125262 341778 125294 342334
rect 123728 331174 124048 331206
rect 123728 330938 123770 331174
rect 124006 330938 124048 331174
rect 123728 330854 124048 330938
rect 123728 330618 123770 330854
rect 124006 330618 124048 330854
rect 123728 330586 124048 330618
rect 120954 302058 120986 302614
rect 121542 302058 121574 302614
rect 120954 266614 121574 302058
rect 124674 306334 125294 341778
rect 124674 305778 124706 306334
rect 125262 305778 125294 306334
rect 123728 295174 124048 295206
rect 123728 294938 123770 295174
rect 124006 294938 124048 295174
rect 123728 294854 124048 294938
rect 123728 294618 123770 294854
rect 124006 294618 124048 294854
rect 123728 294586 124048 294618
rect 120954 266058 120986 266614
rect 121542 266058 121574 266614
rect 120954 230614 121574 266058
rect 124674 270334 125294 305778
rect 124674 269778 124706 270334
rect 125262 269778 125294 270334
rect 123728 259174 124048 259206
rect 123728 258938 123770 259174
rect 124006 258938 124048 259174
rect 123728 258854 124048 258938
rect 123728 258618 123770 258854
rect 124006 258618 124048 258854
rect 123728 258586 124048 258618
rect 120954 230058 120986 230614
rect 121542 230058 121574 230614
rect 120954 194614 121574 230058
rect 124674 234334 125294 269778
rect 124674 233778 124706 234334
rect 125262 233778 125294 234334
rect 123728 223174 124048 223206
rect 123728 222938 123770 223174
rect 124006 222938 124048 223174
rect 123728 222854 124048 222938
rect 123728 222618 123770 222854
rect 124006 222618 124048 222854
rect 123728 222586 124048 222618
rect 120954 194058 120986 194614
rect 121542 194058 121574 194614
rect 120954 158614 121574 194058
rect 124674 198334 125294 233778
rect 124674 197778 124706 198334
rect 125262 197778 125294 198334
rect 123728 187174 124048 187206
rect 123728 186938 123770 187174
rect 124006 186938 124048 187174
rect 123728 186854 124048 186938
rect 123728 186618 123770 186854
rect 124006 186618 124048 186854
rect 123728 186586 124048 186618
rect 120954 158058 120986 158614
rect 121542 158058 121574 158614
rect 120954 122614 121574 158058
rect 124674 162334 125294 197778
rect 124674 161778 124706 162334
rect 125262 161778 125294 162334
rect 123728 151174 124048 151206
rect 123728 150938 123770 151174
rect 124006 150938 124048 151174
rect 123728 150854 124048 150938
rect 123728 150618 123770 150854
rect 124006 150618 124048 150854
rect 123728 150586 124048 150618
rect 120954 122058 120986 122614
rect 121542 122058 121574 122614
rect 120954 86614 121574 122058
rect 124674 126334 125294 161778
rect 124674 125778 124706 126334
rect 125262 125778 125294 126334
rect 123728 115174 124048 115206
rect 123728 114938 123770 115174
rect 124006 114938 124048 115174
rect 123728 114854 124048 114938
rect 123728 114618 123770 114854
rect 124006 114618 124048 114854
rect 123728 114586 124048 114618
rect 120954 86058 120986 86614
rect 121542 86058 121574 86614
rect 120954 50614 121574 86058
rect 124674 90334 125294 125778
rect 124674 89778 124706 90334
rect 125262 89778 125294 90334
rect 123728 79174 124048 79206
rect 123728 78938 123770 79174
rect 124006 78938 124048 79174
rect 123728 78854 124048 78938
rect 123728 78618 123770 78854
rect 124006 78618 124048 78854
rect 123728 78586 124048 78618
rect 120954 50058 120986 50614
rect 121542 50058 121574 50614
rect 120954 14614 121574 50058
rect 124674 54334 125294 89778
rect 124674 53778 124706 54334
rect 125262 53778 125294 54334
rect 123728 43174 124048 43206
rect 123728 42938 123770 43174
rect 124006 42938 124048 43174
rect 123728 42854 124048 42938
rect 123728 42618 123770 42854
rect 124006 42618 124048 42854
rect 123728 42586 124048 42618
rect 120954 14058 120986 14614
rect 121542 14058 121574 14614
rect 120954 -3226 121574 14058
rect 124674 18334 125294 53778
rect 124674 17778 124706 18334
rect 125262 17778 125294 18334
rect 123728 7174 124048 7206
rect 123728 6938 123770 7174
rect 124006 6938 124048 7174
rect 123728 6854 124048 6938
rect 123728 6618 123770 6854
rect 124006 6618 124048 6854
rect 123728 6586 124048 6618
rect 120954 -3782 120986 -3226
rect 121542 -3782 121574 -3226
rect 120954 -7654 121574 -3782
rect 124674 -4186 125294 17778
rect 124674 -4742 124706 -4186
rect 125262 -4742 125294 -4186
rect 124674 -7654 125294 -4742
rect 128394 709638 129014 711590
rect 128394 709082 128426 709638
rect 128982 709082 129014 709638
rect 128394 670054 129014 709082
rect 128394 669498 128426 670054
rect 128982 669498 129014 670054
rect 128394 634054 129014 669498
rect 128394 633498 128426 634054
rect 128982 633498 129014 634054
rect 128394 598054 129014 633498
rect 128394 597498 128426 598054
rect 128982 597498 129014 598054
rect 128394 562054 129014 597498
rect 128394 561498 128426 562054
rect 128982 561498 129014 562054
rect 128394 526054 129014 561498
rect 128394 525498 128426 526054
rect 128982 525498 129014 526054
rect 128394 490054 129014 525498
rect 128394 489498 128426 490054
rect 128982 489498 129014 490054
rect 128394 454054 129014 489498
rect 128394 453498 128426 454054
rect 128982 453498 129014 454054
rect 128394 418054 129014 453498
rect 128394 417498 128426 418054
rect 128982 417498 129014 418054
rect 128394 382054 129014 417498
rect 128394 381498 128426 382054
rect 128982 381498 129014 382054
rect 128394 346054 129014 381498
rect 128394 345498 128426 346054
rect 128982 345498 129014 346054
rect 128394 310054 129014 345498
rect 128394 309498 128426 310054
rect 128982 309498 129014 310054
rect 128394 274054 129014 309498
rect 128394 273498 128426 274054
rect 128982 273498 129014 274054
rect 128394 238054 129014 273498
rect 128394 237498 128426 238054
rect 128982 237498 129014 238054
rect 128394 202054 129014 237498
rect 128394 201498 128426 202054
rect 128982 201498 129014 202054
rect 128394 166054 129014 201498
rect 128394 165498 128426 166054
rect 128982 165498 129014 166054
rect 128394 130054 129014 165498
rect 128394 129498 128426 130054
rect 128982 129498 129014 130054
rect 128394 94054 129014 129498
rect 128394 93498 128426 94054
rect 128982 93498 129014 94054
rect 128394 58054 129014 93498
rect 128394 57498 128426 58054
rect 128982 57498 129014 58054
rect 128394 22054 129014 57498
rect 128394 21498 128426 22054
rect 128982 21498 129014 22054
rect 128394 -5146 129014 21498
rect 128394 -5702 128426 -5146
rect 128982 -5702 129014 -5146
rect 128394 -7654 129014 -5702
rect 132114 710598 132734 711590
rect 132114 710042 132146 710598
rect 132702 710042 132734 710598
rect 132114 673774 132734 710042
rect 132114 673218 132146 673774
rect 132702 673218 132734 673774
rect 132114 637774 132734 673218
rect 132114 637218 132146 637774
rect 132702 637218 132734 637774
rect 132114 601774 132734 637218
rect 132114 601218 132146 601774
rect 132702 601218 132734 601774
rect 132114 565774 132734 601218
rect 132114 565218 132146 565774
rect 132702 565218 132734 565774
rect 132114 529774 132734 565218
rect 132114 529218 132146 529774
rect 132702 529218 132734 529774
rect 132114 493774 132734 529218
rect 132114 493218 132146 493774
rect 132702 493218 132734 493774
rect 132114 457774 132734 493218
rect 132114 457218 132146 457774
rect 132702 457218 132734 457774
rect 132114 421774 132734 457218
rect 132114 421218 132146 421774
rect 132702 421218 132734 421774
rect 132114 385774 132734 421218
rect 132114 385218 132146 385774
rect 132702 385218 132734 385774
rect 132114 349774 132734 385218
rect 132114 349218 132146 349774
rect 132702 349218 132734 349774
rect 132114 313774 132734 349218
rect 132114 313218 132146 313774
rect 132702 313218 132734 313774
rect 132114 277774 132734 313218
rect 132114 277218 132146 277774
rect 132702 277218 132734 277774
rect 132114 241774 132734 277218
rect 132114 241218 132146 241774
rect 132702 241218 132734 241774
rect 132114 205774 132734 241218
rect 132114 205218 132146 205774
rect 132702 205218 132734 205774
rect 132114 169774 132734 205218
rect 132114 169218 132146 169774
rect 132702 169218 132734 169774
rect 132114 133774 132734 169218
rect 132114 133218 132146 133774
rect 132702 133218 132734 133774
rect 132114 97774 132734 133218
rect 132114 97218 132146 97774
rect 132702 97218 132734 97774
rect 132114 61774 132734 97218
rect 132114 61218 132146 61774
rect 132702 61218 132734 61774
rect 132114 25774 132734 61218
rect 132114 25218 132146 25774
rect 132702 25218 132734 25774
rect 132114 -6106 132734 25218
rect 132114 -6662 132146 -6106
rect 132702 -6662 132734 -6106
rect 132114 -7654 132734 -6662
rect 135834 711558 136454 711590
rect 135834 711002 135866 711558
rect 136422 711002 136454 711558
rect 135834 677494 136454 711002
rect 135834 676938 135866 677494
rect 136422 676938 136454 677494
rect 135834 641494 136454 676938
rect 135834 640938 135866 641494
rect 136422 640938 136454 641494
rect 135834 605494 136454 640938
rect 135834 604938 135866 605494
rect 136422 604938 136454 605494
rect 135834 569494 136454 604938
rect 135834 568938 135866 569494
rect 136422 568938 136454 569494
rect 135834 533494 136454 568938
rect 135834 532938 135866 533494
rect 136422 532938 136454 533494
rect 135834 497494 136454 532938
rect 135834 496938 135866 497494
rect 136422 496938 136454 497494
rect 135834 461494 136454 496938
rect 135834 460938 135866 461494
rect 136422 460938 136454 461494
rect 135834 425494 136454 460938
rect 135834 424938 135866 425494
rect 136422 424938 136454 425494
rect 135834 389494 136454 424938
rect 135834 388938 135866 389494
rect 136422 388938 136454 389494
rect 135834 353494 136454 388938
rect 135834 352938 135866 353494
rect 136422 352938 136454 353494
rect 135834 317494 136454 352938
rect 145794 704838 146414 711590
rect 145794 704282 145826 704838
rect 146382 704282 146414 704838
rect 145794 687454 146414 704282
rect 145794 686898 145826 687454
rect 146382 686898 146414 687454
rect 145794 651454 146414 686898
rect 145794 650898 145826 651454
rect 146382 650898 146414 651454
rect 145794 615454 146414 650898
rect 145794 614898 145826 615454
rect 146382 614898 146414 615454
rect 145794 579454 146414 614898
rect 145794 578898 145826 579454
rect 146382 578898 146414 579454
rect 145794 543454 146414 578898
rect 145794 542898 145826 543454
rect 146382 542898 146414 543454
rect 145794 507454 146414 542898
rect 145794 506898 145826 507454
rect 146382 506898 146414 507454
rect 145794 471454 146414 506898
rect 145794 470898 145826 471454
rect 146382 470898 146414 471454
rect 145794 435454 146414 470898
rect 145794 434898 145826 435454
rect 146382 434898 146414 435454
rect 145794 399454 146414 434898
rect 145794 398898 145826 399454
rect 146382 398898 146414 399454
rect 145794 363454 146414 398898
rect 145794 362898 145826 363454
rect 146382 362898 146414 363454
rect 139088 327454 139408 327486
rect 139088 327218 139130 327454
rect 139366 327218 139408 327454
rect 139088 327134 139408 327218
rect 139088 326898 139130 327134
rect 139366 326898 139408 327134
rect 139088 326866 139408 326898
rect 145794 327454 146414 362898
rect 145794 326898 145826 327454
rect 146382 326898 146414 327454
rect 135834 316938 135866 317494
rect 136422 316938 136454 317494
rect 135834 281494 136454 316938
rect 139088 291454 139408 291486
rect 139088 291218 139130 291454
rect 139366 291218 139408 291454
rect 139088 291134 139408 291218
rect 139088 290898 139130 291134
rect 139366 290898 139408 291134
rect 139088 290866 139408 290898
rect 145794 291454 146414 326898
rect 145794 290898 145826 291454
rect 146382 290898 146414 291454
rect 135834 280938 135866 281494
rect 136422 280938 136454 281494
rect 135834 245494 136454 280938
rect 139088 255454 139408 255486
rect 139088 255218 139130 255454
rect 139366 255218 139408 255454
rect 139088 255134 139408 255218
rect 139088 254898 139130 255134
rect 139366 254898 139408 255134
rect 139088 254866 139408 254898
rect 145794 255454 146414 290898
rect 145794 254898 145826 255454
rect 146382 254898 146414 255454
rect 135834 244938 135866 245494
rect 136422 244938 136454 245494
rect 135834 209494 136454 244938
rect 139088 219454 139408 219486
rect 139088 219218 139130 219454
rect 139366 219218 139408 219454
rect 139088 219134 139408 219218
rect 139088 218898 139130 219134
rect 139366 218898 139408 219134
rect 139088 218866 139408 218898
rect 145794 219454 146414 254898
rect 145794 218898 145826 219454
rect 146382 218898 146414 219454
rect 135834 208938 135866 209494
rect 136422 208938 136454 209494
rect 135834 173494 136454 208938
rect 139088 183454 139408 183486
rect 139088 183218 139130 183454
rect 139366 183218 139408 183454
rect 139088 183134 139408 183218
rect 139088 182898 139130 183134
rect 139366 182898 139408 183134
rect 139088 182866 139408 182898
rect 145794 183454 146414 218898
rect 145794 182898 145826 183454
rect 146382 182898 146414 183454
rect 135834 172938 135866 173494
rect 136422 172938 136454 173494
rect 135834 137494 136454 172938
rect 139088 147454 139408 147486
rect 139088 147218 139130 147454
rect 139366 147218 139408 147454
rect 139088 147134 139408 147218
rect 139088 146898 139130 147134
rect 139366 146898 139408 147134
rect 139088 146866 139408 146898
rect 145794 147454 146414 182898
rect 145794 146898 145826 147454
rect 146382 146898 146414 147454
rect 135834 136938 135866 137494
rect 136422 136938 136454 137494
rect 135834 101494 136454 136938
rect 139088 111454 139408 111486
rect 139088 111218 139130 111454
rect 139366 111218 139408 111454
rect 139088 111134 139408 111218
rect 139088 110898 139130 111134
rect 139366 110898 139408 111134
rect 139088 110866 139408 110898
rect 145794 111454 146414 146898
rect 145794 110898 145826 111454
rect 146382 110898 146414 111454
rect 135834 100938 135866 101494
rect 136422 100938 136454 101494
rect 135834 65494 136454 100938
rect 139088 75454 139408 75486
rect 139088 75218 139130 75454
rect 139366 75218 139408 75454
rect 139088 75134 139408 75218
rect 139088 74898 139130 75134
rect 139366 74898 139408 75134
rect 139088 74866 139408 74898
rect 145794 75454 146414 110898
rect 145794 74898 145826 75454
rect 146382 74898 146414 75454
rect 135834 64938 135866 65494
rect 136422 64938 136454 65494
rect 135834 29494 136454 64938
rect 139088 39454 139408 39486
rect 139088 39218 139130 39454
rect 139366 39218 139408 39454
rect 139088 39134 139408 39218
rect 139088 38898 139130 39134
rect 139366 38898 139408 39134
rect 139088 38866 139408 38898
rect 145794 39454 146414 74898
rect 145794 38898 145826 39454
rect 146382 38898 146414 39454
rect 135834 28938 135866 29494
rect 136422 28938 136454 29494
rect 135834 -7066 136454 28938
rect 135834 -7622 135866 -7066
rect 136422 -7622 136454 -7066
rect 135834 -7654 136454 -7622
rect 145794 3454 146414 38898
rect 145794 2898 145826 3454
rect 146382 2898 146414 3454
rect 145794 -346 146414 2898
rect 145794 -902 145826 -346
rect 146382 -902 146414 -346
rect 145794 -7654 146414 -902
rect 149514 705798 150134 711590
rect 149514 705242 149546 705798
rect 150102 705242 150134 705798
rect 149514 691174 150134 705242
rect 149514 690618 149546 691174
rect 150102 690618 150134 691174
rect 149514 655174 150134 690618
rect 149514 654618 149546 655174
rect 150102 654618 150134 655174
rect 149514 619174 150134 654618
rect 149514 618618 149546 619174
rect 150102 618618 150134 619174
rect 149514 583174 150134 618618
rect 149514 582618 149546 583174
rect 150102 582618 150134 583174
rect 149514 547174 150134 582618
rect 149514 546618 149546 547174
rect 150102 546618 150134 547174
rect 149514 511174 150134 546618
rect 149514 510618 149546 511174
rect 150102 510618 150134 511174
rect 149514 475174 150134 510618
rect 149514 474618 149546 475174
rect 150102 474618 150134 475174
rect 149514 439174 150134 474618
rect 149514 438618 149546 439174
rect 150102 438618 150134 439174
rect 149514 403174 150134 438618
rect 149514 402618 149546 403174
rect 150102 402618 150134 403174
rect 149514 367174 150134 402618
rect 149514 366618 149546 367174
rect 150102 366618 150134 367174
rect 149514 331174 150134 366618
rect 149514 330618 149546 331174
rect 150102 330618 150134 331174
rect 149514 295174 150134 330618
rect 149514 294618 149546 295174
rect 150102 294618 150134 295174
rect 149514 259174 150134 294618
rect 149514 258618 149546 259174
rect 150102 258618 150134 259174
rect 149514 223174 150134 258618
rect 149514 222618 149546 223174
rect 150102 222618 150134 223174
rect 149514 187174 150134 222618
rect 149514 186618 149546 187174
rect 150102 186618 150134 187174
rect 149514 151174 150134 186618
rect 149514 150618 149546 151174
rect 150102 150618 150134 151174
rect 149514 115174 150134 150618
rect 149514 114618 149546 115174
rect 150102 114618 150134 115174
rect 149514 79174 150134 114618
rect 149514 78618 149546 79174
rect 150102 78618 150134 79174
rect 149514 43174 150134 78618
rect 149514 42618 149546 43174
rect 150102 42618 150134 43174
rect 149514 7174 150134 42618
rect 149514 6618 149546 7174
rect 150102 6618 150134 7174
rect 149514 -1306 150134 6618
rect 149514 -1862 149546 -1306
rect 150102 -1862 150134 -1306
rect 149514 -7654 150134 -1862
rect 153234 706758 153854 711590
rect 153234 706202 153266 706758
rect 153822 706202 153854 706758
rect 153234 694894 153854 706202
rect 153234 694338 153266 694894
rect 153822 694338 153854 694894
rect 153234 658894 153854 694338
rect 153234 658338 153266 658894
rect 153822 658338 153854 658894
rect 153234 622894 153854 658338
rect 153234 622338 153266 622894
rect 153822 622338 153854 622894
rect 153234 586894 153854 622338
rect 153234 586338 153266 586894
rect 153822 586338 153854 586894
rect 153234 550894 153854 586338
rect 153234 550338 153266 550894
rect 153822 550338 153854 550894
rect 153234 514894 153854 550338
rect 153234 514338 153266 514894
rect 153822 514338 153854 514894
rect 153234 478894 153854 514338
rect 153234 478338 153266 478894
rect 153822 478338 153854 478894
rect 153234 442894 153854 478338
rect 153234 442338 153266 442894
rect 153822 442338 153854 442894
rect 153234 406894 153854 442338
rect 153234 406338 153266 406894
rect 153822 406338 153854 406894
rect 153234 370894 153854 406338
rect 153234 370338 153266 370894
rect 153822 370338 153854 370894
rect 153234 334894 153854 370338
rect 153234 334338 153266 334894
rect 153822 334338 153854 334894
rect 153234 298894 153854 334338
rect 156954 707718 157574 711590
rect 156954 707162 156986 707718
rect 157542 707162 157574 707718
rect 156954 698614 157574 707162
rect 156954 698058 156986 698614
rect 157542 698058 157574 698614
rect 156954 662614 157574 698058
rect 156954 662058 156986 662614
rect 157542 662058 157574 662614
rect 156954 626614 157574 662058
rect 156954 626058 156986 626614
rect 157542 626058 157574 626614
rect 156954 590614 157574 626058
rect 156954 590058 156986 590614
rect 157542 590058 157574 590614
rect 156954 554614 157574 590058
rect 156954 554058 156986 554614
rect 157542 554058 157574 554614
rect 156954 518614 157574 554058
rect 156954 518058 156986 518614
rect 157542 518058 157574 518614
rect 156954 482614 157574 518058
rect 156954 482058 156986 482614
rect 157542 482058 157574 482614
rect 156954 446614 157574 482058
rect 156954 446058 156986 446614
rect 157542 446058 157574 446614
rect 156954 410614 157574 446058
rect 156954 410058 156986 410614
rect 157542 410058 157574 410614
rect 156954 374614 157574 410058
rect 156954 374058 156986 374614
rect 157542 374058 157574 374614
rect 156954 338614 157574 374058
rect 156954 338058 156986 338614
rect 157542 338058 157574 338614
rect 154448 331174 154768 331206
rect 154448 330938 154490 331174
rect 154726 330938 154768 331174
rect 154448 330854 154768 330938
rect 154448 330618 154490 330854
rect 154726 330618 154768 330854
rect 154448 330586 154768 330618
rect 153234 298338 153266 298894
rect 153822 298338 153854 298894
rect 153234 262894 153854 298338
rect 156954 302614 157574 338058
rect 156954 302058 156986 302614
rect 157542 302058 157574 302614
rect 154448 295174 154768 295206
rect 154448 294938 154490 295174
rect 154726 294938 154768 295174
rect 154448 294854 154768 294938
rect 154448 294618 154490 294854
rect 154726 294618 154768 294854
rect 154448 294586 154768 294618
rect 153234 262338 153266 262894
rect 153822 262338 153854 262894
rect 153234 226894 153854 262338
rect 156954 266614 157574 302058
rect 156954 266058 156986 266614
rect 157542 266058 157574 266614
rect 154448 259174 154768 259206
rect 154448 258938 154490 259174
rect 154726 258938 154768 259174
rect 154448 258854 154768 258938
rect 154448 258618 154490 258854
rect 154726 258618 154768 258854
rect 154448 258586 154768 258618
rect 153234 226338 153266 226894
rect 153822 226338 153854 226894
rect 153234 190894 153854 226338
rect 156954 230614 157574 266058
rect 156954 230058 156986 230614
rect 157542 230058 157574 230614
rect 154448 223174 154768 223206
rect 154448 222938 154490 223174
rect 154726 222938 154768 223174
rect 154448 222854 154768 222938
rect 154448 222618 154490 222854
rect 154726 222618 154768 222854
rect 154448 222586 154768 222618
rect 153234 190338 153266 190894
rect 153822 190338 153854 190894
rect 153234 154894 153854 190338
rect 156954 194614 157574 230058
rect 156954 194058 156986 194614
rect 157542 194058 157574 194614
rect 154448 187174 154768 187206
rect 154448 186938 154490 187174
rect 154726 186938 154768 187174
rect 154448 186854 154768 186938
rect 154448 186618 154490 186854
rect 154726 186618 154768 186854
rect 154448 186586 154768 186618
rect 153234 154338 153266 154894
rect 153822 154338 153854 154894
rect 153234 118894 153854 154338
rect 156954 158614 157574 194058
rect 156954 158058 156986 158614
rect 157542 158058 157574 158614
rect 154448 151174 154768 151206
rect 154448 150938 154490 151174
rect 154726 150938 154768 151174
rect 154448 150854 154768 150938
rect 154448 150618 154490 150854
rect 154726 150618 154768 150854
rect 154448 150586 154768 150618
rect 153234 118338 153266 118894
rect 153822 118338 153854 118894
rect 153234 82894 153854 118338
rect 156954 122614 157574 158058
rect 156954 122058 156986 122614
rect 157542 122058 157574 122614
rect 154448 115174 154768 115206
rect 154448 114938 154490 115174
rect 154726 114938 154768 115174
rect 154448 114854 154768 114938
rect 154448 114618 154490 114854
rect 154726 114618 154768 114854
rect 154448 114586 154768 114618
rect 153234 82338 153266 82894
rect 153822 82338 153854 82894
rect 153234 46894 153854 82338
rect 156954 86614 157574 122058
rect 156954 86058 156986 86614
rect 157542 86058 157574 86614
rect 154448 79174 154768 79206
rect 154448 78938 154490 79174
rect 154726 78938 154768 79174
rect 154448 78854 154768 78938
rect 154448 78618 154490 78854
rect 154726 78618 154768 78854
rect 154448 78586 154768 78618
rect 153234 46338 153266 46894
rect 153822 46338 153854 46894
rect 153234 10894 153854 46338
rect 156954 50614 157574 86058
rect 156954 50058 156986 50614
rect 157542 50058 157574 50614
rect 154448 43174 154768 43206
rect 154448 42938 154490 43174
rect 154726 42938 154768 43174
rect 154448 42854 154768 42938
rect 154448 42618 154490 42854
rect 154726 42618 154768 42854
rect 154448 42586 154768 42618
rect 153234 10338 153266 10894
rect 153822 10338 153854 10894
rect 153234 -2266 153854 10338
rect 156954 14614 157574 50058
rect 156954 14058 156986 14614
rect 157542 14058 157574 14614
rect 154448 7174 154768 7206
rect 154448 6938 154490 7174
rect 154726 6938 154768 7174
rect 154448 6854 154768 6938
rect 154448 6618 154490 6854
rect 154726 6618 154768 6854
rect 154448 6586 154768 6618
rect 153234 -2822 153266 -2266
rect 153822 -2822 153854 -2266
rect 153234 -7654 153854 -2822
rect 156954 -3226 157574 14058
rect 156954 -3782 156986 -3226
rect 157542 -3782 157574 -3226
rect 156954 -7654 157574 -3782
rect 160674 708678 161294 711590
rect 160674 708122 160706 708678
rect 161262 708122 161294 708678
rect 160674 666334 161294 708122
rect 160674 665778 160706 666334
rect 161262 665778 161294 666334
rect 160674 630334 161294 665778
rect 160674 629778 160706 630334
rect 161262 629778 161294 630334
rect 160674 594334 161294 629778
rect 160674 593778 160706 594334
rect 161262 593778 161294 594334
rect 160674 558334 161294 593778
rect 160674 557778 160706 558334
rect 161262 557778 161294 558334
rect 160674 522334 161294 557778
rect 160674 521778 160706 522334
rect 161262 521778 161294 522334
rect 160674 486334 161294 521778
rect 160674 485778 160706 486334
rect 161262 485778 161294 486334
rect 160674 450334 161294 485778
rect 160674 449778 160706 450334
rect 161262 449778 161294 450334
rect 160674 414334 161294 449778
rect 160674 413778 160706 414334
rect 161262 413778 161294 414334
rect 160674 378334 161294 413778
rect 160674 377778 160706 378334
rect 161262 377778 161294 378334
rect 160674 342334 161294 377778
rect 160674 341778 160706 342334
rect 161262 341778 161294 342334
rect 160674 306334 161294 341778
rect 160674 305778 160706 306334
rect 161262 305778 161294 306334
rect 160674 270334 161294 305778
rect 160674 269778 160706 270334
rect 161262 269778 161294 270334
rect 160674 234334 161294 269778
rect 160674 233778 160706 234334
rect 161262 233778 161294 234334
rect 160674 198334 161294 233778
rect 160674 197778 160706 198334
rect 161262 197778 161294 198334
rect 160674 162334 161294 197778
rect 160674 161778 160706 162334
rect 161262 161778 161294 162334
rect 160674 126334 161294 161778
rect 160674 125778 160706 126334
rect 161262 125778 161294 126334
rect 160674 90334 161294 125778
rect 160674 89778 160706 90334
rect 161262 89778 161294 90334
rect 160674 54334 161294 89778
rect 160674 53778 160706 54334
rect 161262 53778 161294 54334
rect 160674 18334 161294 53778
rect 160674 17778 160706 18334
rect 161262 17778 161294 18334
rect 160674 -4186 161294 17778
rect 160674 -4742 160706 -4186
rect 161262 -4742 161294 -4186
rect 160674 -7654 161294 -4742
rect 164394 709638 165014 711590
rect 164394 709082 164426 709638
rect 164982 709082 165014 709638
rect 164394 670054 165014 709082
rect 164394 669498 164426 670054
rect 164982 669498 165014 670054
rect 164394 634054 165014 669498
rect 164394 633498 164426 634054
rect 164982 633498 165014 634054
rect 164394 598054 165014 633498
rect 164394 597498 164426 598054
rect 164982 597498 165014 598054
rect 164394 562054 165014 597498
rect 164394 561498 164426 562054
rect 164982 561498 165014 562054
rect 164394 526054 165014 561498
rect 164394 525498 164426 526054
rect 164982 525498 165014 526054
rect 164394 490054 165014 525498
rect 164394 489498 164426 490054
rect 164982 489498 165014 490054
rect 164394 454054 165014 489498
rect 164394 453498 164426 454054
rect 164982 453498 165014 454054
rect 164394 418054 165014 453498
rect 164394 417498 164426 418054
rect 164982 417498 165014 418054
rect 164394 382054 165014 417498
rect 164394 381498 164426 382054
rect 164982 381498 165014 382054
rect 164394 346054 165014 381498
rect 164394 345498 164426 346054
rect 164982 345498 165014 346054
rect 164394 310054 165014 345498
rect 164394 309498 164426 310054
rect 164982 309498 165014 310054
rect 164394 274054 165014 309498
rect 164394 273498 164426 274054
rect 164982 273498 165014 274054
rect 164394 238054 165014 273498
rect 164394 237498 164426 238054
rect 164982 237498 165014 238054
rect 164394 202054 165014 237498
rect 164394 201498 164426 202054
rect 164982 201498 165014 202054
rect 164394 166054 165014 201498
rect 164394 165498 164426 166054
rect 164982 165498 165014 166054
rect 164394 130054 165014 165498
rect 164394 129498 164426 130054
rect 164982 129498 165014 130054
rect 164394 94054 165014 129498
rect 164394 93498 164426 94054
rect 164982 93498 165014 94054
rect 164394 58054 165014 93498
rect 164394 57498 164426 58054
rect 164982 57498 165014 58054
rect 164394 22054 165014 57498
rect 164394 21498 164426 22054
rect 164982 21498 165014 22054
rect 164394 -5146 165014 21498
rect 164394 -5702 164426 -5146
rect 164982 -5702 165014 -5146
rect 164394 -7654 165014 -5702
rect 168114 710598 168734 711590
rect 168114 710042 168146 710598
rect 168702 710042 168734 710598
rect 168114 673774 168734 710042
rect 168114 673218 168146 673774
rect 168702 673218 168734 673774
rect 168114 637774 168734 673218
rect 168114 637218 168146 637774
rect 168702 637218 168734 637774
rect 168114 601774 168734 637218
rect 168114 601218 168146 601774
rect 168702 601218 168734 601774
rect 168114 565774 168734 601218
rect 168114 565218 168146 565774
rect 168702 565218 168734 565774
rect 168114 529774 168734 565218
rect 168114 529218 168146 529774
rect 168702 529218 168734 529774
rect 168114 493774 168734 529218
rect 168114 493218 168146 493774
rect 168702 493218 168734 493774
rect 168114 457774 168734 493218
rect 168114 457218 168146 457774
rect 168702 457218 168734 457774
rect 168114 421774 168734 457218
rect 168114 421218 168146 421774
rect 168702 421218 168734 421774
rect 168114 385774 168734 421218
rect 168114 385218 168146 385774
rect 168702 385218 168734 385774
rect 168114 349774 168734 385218
rect 168114 349218 168146 349774
rect 168702 349218 168734 349774
rect 168114 313774 168734 349218
rect 171834 711558 172454 711590
rect 171834 711002 171866 711558
rect 172422 711002 172454 711558
rect 171834 677494 172454 711002
rect 171834 676938 171866 677494
rect 172422 676938 172454 677494
rect 171834 641494 172454 676938
rect 171834 640938 171866 641494
rect 172422 640938 172454 641494
rect 171834 605494 172454 640938
rect 171834 604938 171866 605494
rect 172422 604938 172454 605494
rect 171834 569494 172454 604938
rect 171834 568938 171866 569494
rect 172422 568938 172454 569494
rect 171834 533494 172454 568938
rect 171834 532938 171866 533494
rect 172422 532938 172454 533494
rect 171834 497494 172454 532938
rect 171834 496938 171866 497494
rect 172422 496938 172454 497494
rect 171834 461494 172454 496938
rect 171834 460938 171866 461494
rect 172422 460938 172454 461494
rect 171834 425494 172454 460938
rect 171834 424938 171866 425494
rect 172422 424938 172454 425494
rect 171834 389494 172454 424938
rect 171834 388938 171866 389494
rect 172422 388938 172454 389494
rect 171834 353494 172454 388938
rect 171834 352938 171866 353494
rect 172422 352938 172454 353494
rect 169808 327454 170128 327486
rect 169808 327218 169850 327454
rect 170086 327218 170128 327454
rect 169808 327134 170128 327218
rect 169808 326898 169850 327134
rect 170086 326898 170128 327134
rect 169808 326866 170128 326898
rect 168114 313218 168146 313774
rect 168702 313218 168734 313774
rect 168114 277774 168734 313218
rect 171834 317494 172454 352938
rect 171834 316938 171866 317494
rect 172422 316938 172454 317494
rect 169808 291454 170128 291486
rect 169808 291218 169850 291454
rect 170086 291218 170128 291454
rect 169808 291134 170128 291218
rect 169808 290898 169850 291134
rect 170086 290898 170128 291134
rect 169808 290866 170128 290898
rect 168114 277218 168146 277774
rect 168702 277218 168734 277774
rect 168114 241774 168734 277218
rect 171834 281494 172454 316938
rect 171834 280938 171866 281494
rect 172422 280938 172454 281494
rect 169808 255454 170128 255486
rect 169808 255218 169850 255454
rect 170086 255218 170128 255454
rect 169808 255134 170128 255218
rect 169808 254898 169850 255134
rect 170086 254898 170128 255134
rect 169808 254866 170128 254898
rect 168114 241218 168146 241774
rect 168702 241218 168734 241774
rect 168114 205774 168734 241218
rect 171834 245494 172454 280938
rect 171834 244938 171866 245494
rect 172422 244938 172454 245494
rect 169808 219454 170128 219486
rect 169808 219218 169850 219454
rect 170086 219218 170128 219454
rect 169808 219134 170128 219218
rect 169808 218898 169850 219134
rect 170086 218898 170128 219134
rect 169808 218866 170128 218898
rect 168114 205218 168146 205774
rect 168702 205218 168734 205774
rect 168114 169774 168734 205218
rect 171834 209494 172454 244938
rect 171834 208938 171866 209494
rect 172422 208938 172454 209494
rect 169808 183454 170128 183486
rect 169808 183218 169850 183454
rect 170086 183218 170128 183454
rect 169808 183134 170128 183218
rect 169808 182898 169850 183134
rect 170086 182898 170128 183134
rect 169808 182866 170128 182898
rect 168114 169218 168146 169774
rect 168702 169218 168734 169774
rect 168114 133774 168734 169218
rect 171834 173494 172454 208938
rect 171834 172938 171866 173494
rect 172422 172938 172454 173494
rect 169808 147454 170128 147486
rect 169808 147218 169850 147454
rect 170086 147218 170128 147454
rect 169808 147134 170128 147218
rect 169808 146898 169850 147134
rect 170086 146898 170128 147134
rect 169808 146866 170128 146898
rect 168114 133218 168146 133774
rect 168702 133218 168734 133774
rect 168114 97774 168734 133218
rect 171834 137494 172454 172938
rect 171834 136938 171866 137494
rect 172422 136938 172454 137494
rect 169808 111454 170128 111486
rect 169808 111218 169850 111454
rect 170086 111218 170128 111454
rect 169808 111134 170128 111218
rect 169808 110898 169850 111134
rect 170086 110898 170128 111134
rect 169808 110866 170128 110898
rect 168114 97218 168146 97774
rect 168702 97218 168734 97774
rect 168114 61774 168734 97218
rect 171834 101494 172454 136938
rect 171834 100938 171866 101494
rect 172422 100938 172454 101494
rect 169808 75454 170128 75486
rect 169808 75218 169850 75454
rect 170086 75218 170128 75454
rect 169808 75134 170128 75218
rect 169808 74898 169850 75134
rect 170086 74898 170128 75134
rect 169808 74866 170128 74898
rect 168114 61218 168146 61774
rect 168702 61218 168734 61774
rect 168114 25774 168734 61218
rect 171834 65494 172454 100938
rect 171834 64938 171866 65494
rect 172422 64938 172454 65494
rect 169808 39454 170128 39486
rect 169808 39218 169850 39454
rect 170086 39218 170128 39454
rect 169808 39134 170128 39218
rect 169808 38898 169850 39134
rect 170086 38898 170128 39134
rect 169808 38866 170128 38898
rect 168114 25218 168146 25774
rect 168702 25218 168734 25774
rect 168114 -6106 168734 25218
rect 168114 -6662 168146 -6106
rect 168702 -6662 168734 -6106
rect 168114 -7654 168734 -6662
rect 171834 29494 172454 64938
rect 171834 28938 171866 29494
rect 172422 28938 172454 29494
rect 171834 -7066 172454 28938
rect 171834 -7622 171866 -7066
rect 172422 -7622 172454 -7066
rect 171834 -7654 172454 -7622
rect 181794 704838 182414 711590
rect 181794 704282 181826 704838
rect 182382 704282 182414 704838
rect 181794 687454 182414 704282
rect 181794 686898 181826 687454
rect 182382 686898 182414 687454
rect 181794 651454 182414 686898
rect 181794 650898 181826 651454
rect 182382 650898 182414 651454
rect 181794 615454 182414 650898
rect 181794 614898 181826 615454
rect 182382 614898 182414 615454
rect 181794 579454 182414 614898
rect 181794 578898 181826 579454
rect 182382 578898 182414 579454
rect 181794 543454 182414 578898
rect 181794 542898 181826 543454
rect 182382 542898 182414 543454
rect 181794 507454 182414 542898
rect 181794 506898 181826 507454
rect 182382 506898 182414 507454
rect 181794 471454 182414 506898
rect 181794 470898 181826 471454
rect 182382 470898 182414 471454
rect 181794 435454 182414 470898
rect 181794 434898 181826 435454
rect 182382 434898 182414 435454
rect 181794 399454 182414 434898
rect 181794 398898 181826 399454
rect 182382 398898 182414 399454
rect 181794 363454 182414 398898
rect 181794 362898 181826 363454
rect 182382 362898 182414 363454
rect 181794 327454 182414 362898
rect 185514 705798 186134 711590
rect 185514 705242 185546 705798
rect 186102 705242 186134 705798
rect 185514 691174 186134 705242
rect 185514 690618 185546 691174
rect 186102 690618 186134 691174
rect 185514 655174 186134 690618
rect 185514 654618 185546 655174
rect 186102 654618 186134 655174
rect 185514 619174 186134 654618
rect 185514 618618 185546 619174
rect 186102 618618 186134 619174
rect 185514 583174 186134 618618
rect 185514 582618 185546 583174
rect 186102 582618 186134 583174
rect 185514 547174 186134 582618
rect 185514 546618 185546 547174
rect 186102 546618 186134 547174
rect 185514 511174 186134 546618
rect 185514 510618 185546 511174
rect 186102 510618 186134 511174
rect 185514 475174 186134 510618
rect 185514 474618 185546 475174
rect 186102 474618 186134 475174
rect 185514 439174 186134 474618
rect 185514 438618 185546 439174
rect 186102 438618 186134 439174
rect 185514 403174 186134 438618
rect 185514 402618 185546 403174
rect 186102 402618 186134 403174
rect 185514 367174 186134 402618
rect 185514 366618 185546 367174
rect 186102 366618 186134 367174
rect 185514 354900 186134 366618
rect 189234 706758 189854 711590
rect 189234 706202 189266 706758
rect 189822 706202 189854 706758
rect 189234 694894 189854 706202
rect 189234 694338 189266 694894
rect 189822 694338 189854 694894
rect 189234 658894 189854 694338
rect 189234 658338 189266 658894
rect 189822 658338 189854 658894
rect 189234 622894 189854 658338
rect 189234 622338 189266 622894
rect 189822 622338 189854 622894
rect 189234 586894 189854 622338
rect 189234 586338 189266 586894
rect 189822 586338 189854 586894
rect 189234 550894 189854 586338
rect 189234 550338 189266 550894
rect 189822 550338 189854 550894
rect 189234 514894 189854 550338
rect 189234 514338 189266 514894
rect 189822 514338 189854 514894
rect 189234 478894 189854 514338
rect 189234 478338 189266 478894
rect 189822 478338 189854 478894
rect 189234 442894 189854 478338
rect 189234 442338 189266 442894
rect 189822 442338 189854 442894
rect 189234 406894 189854 442338
rect 189234 406338 189266 406894
rect 189822 406338 189854 406894
rect 189234 370894 189854 406338
rect 189234 370338 189266 370894
rect 189822 370338 189854 370894
rect 189234 334894 189854 370338
rect 189234 334338 189266 334894
rect 189822 334338 189854 334894
rect 185168 331174 185488 331206
rect 185168 330938 185210 331174
rect 185446 330938 185488 331174
rect 185168 330854 185488 330938
rect 185168 330618 185210 330854
rect 185446 330618 185488 330854
rect 185168 330586 185488 330618
rect 181794 326898 181826 327454
rect 182382 326898 182414 327454
rect 181794 291454 182414 326898
rect 189234 298894 189854 334338
rect 189234 298338 189266 298894
rect 189822 298338 189854 298894
rect 185168 295174 185488 295206
rect 185168 294938 185210 295174
rect 185446 294938 185488 295174
rect 185168 294854 185488 294938
rect 185168 294618 185210 294854
rect 185446 294618 185488 294854
rect 185168 294586 185488 294618
rect 181794 290898 181826 291454
rect 182382 290898 182414 291454
rect 181794 255454 182414 290898
rect 189234 262894 189854 298338
rect 189234 262338 189266 262894
rect 189822 262338 189854 262894
rect 185168 259174 185488 259206
rect 185168 258938 185210 259174
rect 185446 258938 185488 259174
rect 185168 258854 185488 258938
rect 185168 258618 185210 258854
rect 185446 258618 185488 258854
rect 185168 258586 185488 258618
rect 181794 254898 181826 255454
rect 182382 254898 182414 255454
rect 181794 219454 182414 254898
rect 189234 226894 189854 262338
rect 189234 226338 189266 226894
rect 189822 226338 189854 226894
rect 185168 223174 185488 223206
rect 185168 222938 185210 223174
rect 185446 222938 185488 223174
rect 185168 222854 185488 222938
rect 185168 222618 185210 222854
rect 185446 222618 185488 222854
rect 185168 222586 185488 222618
rect 181794 218898 181826 219454
rect 182382 218898 182414 219454
rect 181794 183454 182414 218898
rect 189234 190894 189854 226338
rect 189234 190338 189266 190894
rect 189822 190338 189854 190894
rect 185168 187174 185488 187206
rect 185168 186938 185210 187174
rect 185446 186938 185488 187174
rect 185168 186854 185488 186938
rect 185168 186618 185210 186854
rect 185446 186618 185488 186854
rect 185168 186586 185488 186618
rect 181794 182898 181826 183454
rect 182382 182898 182414 183454
rect 181794 147454 182414 182898
rect 189234 154894 189854 190338
rect 189234 154338 189266 154894
rect 189822 154338 189854 154894
rect 185168 151174 185488 151206
rect 185168 150938 185210 151174
rect 185446 150938 185488 151174
rect 185168 150854 185488 150938
rect 185168 150618 185210 150854
rect 185446 150618 185488 150854
rect 185168 150586 185488 150618
rect 181794 146898 181826 147454
rect 182382 146898 182414 147454
rect 181794 111454 182414 146898
rect 189234 118894 189854 154338
rect 189234 118338 189266 118894
rect 189822 118338 189854 118894
rect 185168 115174 185488 115206
rect 185168 114938 185210 115174
rect 185446 114938 185488 115174
rect 185168 114854 185488 114938
rect 185168 114618 185210 114854
rect 185446 114618 185488 114854
rect 185168 114586 185488 114618
rect 181794 110898 181826 111454
rect 182382 110898 182414 111454
rect 181794 75454 182414 110898
rect 189234 82894 189854 118338
rect 189234 82338 189266 82894
rect 189822 82338 189854 82894
rect 185168 79174 185488 79206
rect 185168 78938 185210 79174
rect 185446 78938 185488 79174
rect 185168 78854 185488 78938
rect 185168 78618 185210 78854
rect 185446 78618 185488 78854
rect 185168 78586 185488 78618
rect 181794 74898 181826 75454
rect 182382 74898 182414 75454
rect 181794 39454 182414 74898
rect 189234 46894 189854 82338
rect 189234 46338 189266 46894
rect 189822 46338 189854 46894
rect 185168 43174 185488 43206
rect 185168 42938 185210 43174
rect 185446 42938 185488 43174
rect 185168 42854 185488 42938
rect 185168 42618 185210 42854
rect 185446 42618 185488 42854
rect 185168 42586 185488 42618
rect 181794 38898 181826 39454
rect 182382 38898 182414 39454
rect 181794 3454 182414 38898
rect 189234 10894 189854 46338
rect 189234 10338 189266 10894
rect 189822 10338 189854 10894
rect 185168 7174 185488 7206
rect 185168 6938 185210 7174
rect 185446 6938 185488 7174
rect 185168 6854 185488 6938
rect 185168 6618 185210 6854
rect 185446 6618 185488 6854
rect 185168 6586 185488 6618
rect 181794 2898 181826 3454
rect 182382 2898 182414 3454
rect 181794 -346 182414 2898
rect 181794 -902 181826 -346
rect 182382 -902 182414 -346
rect 181794 -7654 182414 -902
rect 189234 -2266 189854 10338
rect 189234 -2822 189266 -2266
rect 189822 -2822 189854 -2266
rect 189234 -7654 189854 -2822
rect 192954 707718 193574 711590
rect 192954 707162 192986 707718
rect 193542 707162 193574 707718
rect 192954 698614 193574 707162
rect 192954 698058 192986 698614
rect 193542 698058 193574 698614
rect 192954 662614 193574 698058
rect 192954 662058 192986 662614
rect 193542 662058 193574 662614
rect 192954 626614 193574 662058
rect 192954 626058 192986 626614
rect 193542 626058 193574 626614
rect 192954 590614 193574 626058
rect 192954 590058 192986 590614
rect 193542 590058 193574 590614
rect 192954 554614 193574 590058
rect 192954 554058 192986 554614
rect 193542 554058 193574 554614
rect 192954 518614 193574 554058
rect 192954 518058 192986 518614
rect 193542 518058 193574 518614
rect 192954 482614 193574 518058
rect 192954 482058 192986 482614
rect 193542 482058 193574 482614
rect 192954 446614 193574 482058
rect 192954 446058 192986 446614
rect 193542 446058 193574 446614
rect 192954 410614 193574 446058
rect 192954 410058 192986 410614
rect 193542 410058 193574 410614
rect 192954 374614 193574 410058
rect 192954 374058 192986 374614
rect 193542 374058 193574 374614
rect 192954 338614 193574 374058
rect 192954 338058 192986 338614
rect 193542 338058 193574 338614
rect 192954 302614 193574 338058
rect 192954 302058 192986 302614
rect 193542 302058 193574 302614
rect 192954 266614 193574 302058
rect 192954 266058 192986 266614
rect 193542 266058 193574 266614
rect 192954 230614 193574 266058
rect 192954 230058 192986 230614
rect 193542 230058 193574 230614
rect 192954 194614 193574 230058
rect 192954 194058 192986 194614
rect 193542 194058 193574 194614
rect 192954 158614 193574 194058
rect 192954 158058 192986 158614
rect 193542 158058 193574 158614
rect 192954 122614 193574 158058
rect 192954 122058 192986 122614
rect 193542 122058 193574 122614
rect 192954 86614 193574 122058
rect 192954 86058 192986 86614
rect 193542 86058 193574 86614
rect 192954 50614 193574 86058
rect 192954 50058 192986 50614
rect 193542 50058 193574 50614
rect 192954 14614 193574 50058
rect 192954 14058 192986 14614
rect 193542 14058 193574 14614
rect 192954 -3226 193574 14058
rect 192954 -3782 192986 -3226
rect 193542 -3782 193574 -3226
rect 192954 -7654 193574 -3782
rect 196674 708678 197294 711590
rect 196674 708122 196706 708678
rect 197262 708122 197294 708678
rect 196674 666334 197294 708122
rect 196674 665778 196706 666334
rect 197262 665778 197294 666334
rect 196674 630334 197294 665778
rect 196674 629778 196706 630334
rect 197262 629778 197294 630334
rect 196674 594334 197294 629778
rect 196674 593778 196706 594334
rect 197262 593778 197294 594334
rect 196674 558334 197294 593778
rect 196674 557778 196706 558334
rect 197262 557778 197294 558334
rect 196674 522334 197294 557778
rect 196674 521778 196706 522334
rect 197262 521778 197294 522334
rect 196674 486334 197294 521778
rect 196674 485778 196706 486334
rect 197262 485778 197294 486334
rect 196674 450334 197294 485778
rect 196674 449778 196706 450334
rect 197262 449778 197294 450334
rect 196674 414334 197294 449778
rect 196674 413778 196706 414334
rect 197262 413778 197294 414334
rect 196674 378334 197294 413778
rect 196674 377778 196706 378334
rect 197262 377778 197294 378334
rect 196674 342334 197294 377778
rect 200394 709638 201014 711590
rect 200394 709082 200426 709638
rect 200982 709082 201014 709638
rect 200394 670054 201014 709082
rect 200394 669498 200426 670054
rect 200982 669498 201014 670054
rect 200394 634054 201014 669498
rect 200394 633498 200426 634054
rect 200982 633498 201014 634054
rect 200394 598054 201014 633498
rect 200394 597498 200426 598054
rect 200982 597498 201014 598054
rect 200394 562054 201014 597498
rect 200394 561498 200426 562054
rect 200982 561498 201014 562054
rect 200394 526054 201014 561498
rect 200394 525498 200426 526054
rect 200982 525498 201014 526054
rect 200394 490054 201014 525498
rect 200394 489498 200426 490054
rect 200982 489498 201014 490054
rect 200394 454054 201014 489498
rect 200394 453498 200426 454054
rect 200982 453498 201014 454054
rect 200394 418054 201014 453498
rect 200394 417498 200426 418054
rect 200982 417498 201014 418054
rect 200394 382054 201014 417498
rect 200394 381498 200426 382054
rect 200982 381498 201014 382054
rect 200394 354900 201014 381498
rect 204114 710598 204734 711590
rect 204114 710042 204146 710598
rect 204702 710042 204734 710598
rect 204114 673774 204734 710042
rect 204114 673218 204146 673774
rect 204702 673218 204734 673774
rect 204114 637774 204734 673218
rect 204114 637218 204146 637774
rect 204702 637218 204734 637774
rect 204114 601774 204734 637218
rect 204114 601218 204146 601774
rect 204702 601218 204734 601774
rect 204114 565774 204734 601218
rect 204114 565218 204146 565774
rect 204702 565218 204734 565774
rect 204114 529774 204734 565218
rect 204114 529218 204146 529774
rect 204702 529218 204734 529774
rect 204114 493774 204734 529218
rect 204114 493218 204146 493774
rect 204702 493218 204734 493774
rect 204114 457774 204734 493218
rect 204114 457218 204146 457774
rect 204702 457218 204734 457774
rect 204114 421774 204734 457218
rect 204114 421218 204146 421774
rect 204702 421218 204734 421774
rect 204114 385774 204734 421218
rect 204114 385218 204146 385774
rect 204702 385218 204734 385774
rect 196674 341778 196706 342334
rect 197262 341778 197294 342334
rect 196674 306334 197294 341778
rect 204114 349774 204734 385218
rect 204114 349218 204146 349774
rect 204702 349218 204734 349774
rect 200528 327454 200848 327486
rect 200528 327218 200570 327454
rect 200806 327218 200848 327454
rect 200528 327134 200848 327218
rect 200528 326898 200570 327134
rect 200806 326898 200848 327134
rect 200528 326866 200848 326898
rect 196674 305778 196706 306334
rect 197262 305778 197294 306334
rect 196674 270334 197294 305778
rect 204114 313774 204734 349218
rect 204114 313218 204146 313774
rect 204702 313218 204734 313774
rect 200528 291454 200848 291486
rect 200528 291218 200570 291454
rect 200806 291218 200848 291454
rect 200528 291134 200848 291218
rect 200528 290898 200570 291134
rect 200806 290898 200848 291134
rect 200528 290866 200848 290898
rect 196674 269778 196706 270334
rect 197262 269778 197294 270334
rect 196674 234334 197294 269778
rect 204114 277774 204734 313218
rect 204114 277218 204146 277774
rect 204702 277218 204734 277774
rect 200528 255454 200848 255486
rect 200528 255218 200570 255454
rect 200806 255218 200848 255454
rect 200528 255134 200848 255218
rect 200528 254898 200570 255134
rect 200806 254898 200848 255134
rect 200528 254866 200848 254898
rect 196674 233778 196706 234334
rect 197262 233778 197294 234334
rect 196674 198334 197294 233778
rect 204114 241774 204734 277218
rect 204114 241218 204146 241774
rect 204702 241218 204734 241774
rect 200528 219454 200848 219486
rect 200528 219218 200570 219454
rect 200806 219218 200848 219454
rect 200528 219134 200848 219218
rect 200528 218898 200570 219134
rect 200806 218898 200848 219134
rect 200528 218866 200848 218898
rect 196674 197778 196706 198334
rect 197262 197778 197294 198334
rect 196674 162334 197294 197778
rect 204114 205774 204734 241218
rect 204114 205218 204146 205774
rect 204702 205218 204734 205774
rect 200528 183454 200848 183486
rect 200528 183218 200570 183454
rect 200806 183218 200848 183454
rect 200528 183134 200848 183218
rect 200528 182898 200570 183134
rect 200806 182898 200848 183134
rect 200528 182866 200848 182898
rect 196674 161778 196706 162334
rect 197262 161778 197294 162334
rect 196674 126334 197294 161778
rect 204114 169774 204734 205218
rect 204114 169218 204146 169774
rect 204702 169218 204734 169774
rect 200528 147454 200848 147486
rect 200528 147218 200570 147454
rect 200806 147218 200848 147454
rect 200528 147134 200848 147218
rect 200528 146898 200570 147134
rect 200806 146898 200848 147134
rect 200528 146866 200848 146898
rect 196674 125778 196706 126334
rect 197262 125778 197294 126334
rect 196674 90334 197294 125778
rect 204114 133774 204734 169218
rect 204114 133218 204146 133774
rect 204702 133218 204734 133774
rect 200528 111454 200848 111486
rect 200528 111218 200570 111454
rect 200806 111218 200848 111454
rect 200528 111134 200848 111218
rect 200528 110898 200570 111134
rect 200806 110898 200848 111134
rect 200528 110866 200848 110898
rect 196674 89778 196706 90334
rect 197262 89778 197294 90334
rect 196674 54334 197294 89778
rect 204114 97774 204734 133218
rect 204114 97218 204146 97774
rect 204702 97218 204734 97774
rect 200528 75454 200848 75486
rect 200528 75218 200570 75454
rect 200806 75218 200848 75454
rect 200528 75134 200848 75218
rect 200528 74898 200570 75134
rect 200806 74898 200848 75134
rect 200528 74866 200848 74898
rect 196674 53778 196706 54334
rect 197262 53778 197294 54334
rect 196674 18334 197294 53778
rect 204114 61774 204734 97218
rect 204114 61218 204146 61774
rect 204702 61218 204734 61774
rect 200528 39454 200848 39486
rect 200528 39218 200570 39454
rect 200806 39218 200848 39454
rect 200528 39134 200848 39218
rect 200528 38898 200570 39134
rect 200806 38898 200848 39134
rect 200528 38866 200848 38898
rect 196674 17778 196706 18334
rect 197262 17778 197294 18334
rect 196674 -4186 197294 17778
rect 196674 -4742 196706 -4186
rect 197262 -4742 197294 -4186
rect 196674 -7654 197294 -4742
rect 204114 25774 204734 61218
rect 204114 25218 204146 25774
rect 204702 25218 204734 25774
rect 204114 -6106 204734 25218
rect 204114 -6662 204146 -6106
rect 204702 -6662 204734 -6106
rect 204114 -7654 204734 -6662
rect 207834 711558 208454 711590
rect 207834 711002 207866 711558
rect 208422 711002 208454 711558
rect 207834 677494 208454 711002
rect 207834 676938 207866 677494
rect 208422 676938 208454 677494
rect 207834 641494 208454 676938
rect 207834 640938 207866 641494
rect 208422 640938 208454 641494
rect 207834 605494 208454 640938
rect 207834 604938 207866 605494
rect 208422 604938 208454 605494
rect 207834 569494 208454 604938
rect 207834 568938 207866 569494
rect 208422 568938 208454 569494
rect 207834 533494 208454 568938
rect 207834 532938 207866 533494
rect 208422 532938 208454 533494
rect 207834 497494 208454 532938
rect 207834 496938 207866 497494
rect 208422 496938 208454 497494
rect 207834 461494 208454 496938
rect 207834 460938 207866 461494
rect 208422 460938 208454 461494
rect 207834 425494 208454 460938
rect 207834 424938 207866 425494
rect 208422 424938 208454 425494
rect 207834 389494 208454 424938
rect 207834 388938 207866 389494
rect 208422 388938 208454 389494
rect 207834 353494 208454 388938
rect 207834 352938 207866 353494
rect 208422 352938 208454 353494
rect 207834 317494 208454 352938
rect 217794 704838 218414 711590
rect 217794 704282 217826 704838
rect 218382 704282 218414 704838
rect 217794 687454 218414 704282
rect 217794 686898 217826 687454
rect 218382 686898 218414 687454
rect 217794 651454 218414 686898
rect 217794 650898 217826 651454
rect 218382 650898 218414 651454
rect 217794 615454 218414 650898
rect 217794 614898 217826 615454
rect 218382 614898 218414 615454
rect 217794 579454 218414 614898
rect 217794 578898 217826 579454
rect 218382 578898 218414 579454
rect 217794 543454 218414 578898
rect 217794 542898 217826 543454
rect 218382 542898 218414 543454
rect 217794 507454 218414 542898
rect 217794 506898 217826 507454
rect 218382 506898 218414 507454
rect 217794 471454 218414 506898
rect 217794 470898 217826 471454
rect 218382 470898 218414 471454
rect 217794 435454 218414 470898
rect 217794 434898 217826 435454
rect 218382 434898 218414 435454
rect 217794 399454 218414 434898
rect 217794 398898 217826 399454
rect 218382 398898 218414 399454
rect 217794 363454 218414 398898
rect 217794 362898 217826 363454
rect 218382 362898 218414 363454
rect 215888 331174 216208 331206
rect 215888 330938 215930 331174
rect 216166 330938 216208 331174
rect 215888 330854 216208 330938
rect 215888 330618 215930 330854
rect 216166 330618 216208 330854
rect 215888 330586 216208 330618
rect 207834 316938 207866 317494
rect 208422 316938 208454 317494
rect 207834 281494 208454 316938
rect 217794 327454 218414 362898
rect 217794 326898 217826 327454
rect 218382 326898 218414 327454
rect 215888 295174 216208 295206
rect 215888 294938 215930 295174
rect 216166 294938 216208 295174
rect 215888 294854 216208 294938
rect 215888 294618 215930 294854
rect 216166 294618 216208 294854
rect 215888 294586 216208 294618
rect 207834 280938 207866 281494
rect 208422 280938 208454 281494
rect 207834 245494 208454 280938
rect 217794 291454 218414 326898
rect 217794 290898 217826 291454
rect 218382 290898 218414 291454
rect 215888 259174 216208 259206
rect 215888 258938 215930 259174
rect 216166 258938 216208 259174
rect 215888 258854 216208 258938
rect 215888 258618 215930 258854
rect 216166 258618 216208 258854
rect 215888 258586 216208 258618
rect 207834 244938 207866 245494
rect 208422 244938 208454 245494
rect 207834 209494 208454 244938
rect 217794 255454 218414 290898
rect 217794 254898 217826 255454
rect 218382 254898 218414 255454
rect 215888 223174 216208 223206
rect 215888 222938 215930 223174
rect 216166 222938 216208 223174
rect 215888 222854 216208 222938
rect 215888 222618 215930 222854
rect 216166 222618 216208 222854
rect 215888 222586 216208 222618
rect 207834 208938 207866 209494
rect 208422 208938 208454 209494
rect 207834 173494 208454 208938
rect 217794 219454 218414 254898
rect 217794 218898 217826 219454
rect 218382 218898 218414 219454
rect 215888 187174 216208 187206
rect 215888 186938 215930 187174
rect 216166 186938 216208 187174
rect 215888 186854 216208 186938
rect 215888 186618 215930 186854
rect 216166 186618 216208 186854
rect 215888 186586 216208 186618
rect 207834 172938 207866 173494
rect 208422 172938 208454 173494
rect 207834 137494 208454 172938
rect 217794 183454 218414 218898
rect 217794 182898 217826 183454
rect 218382 182898 218414 183454
rect 215888 151174 216208 151206
rect 215888 150938 215930 151174
rect 216166 150938 216208 151174
rect 215888 150854 216208 150938
rect 215888 150618 215930 150854
rect 216166 150618 216208 150854
rect 215888 150586 216208 150618
rect 207834 136938 207866 137494
rect 208422 136938 208454 137494
rect 207834 101494 208454 136938
rect 217794 147454 218414 182898
rect 217794 146898 217826 147454
rect 218382 146898 218414 147454
rect 215888 115174 216208 115206
rect 215888 114938 215930 115174
rect 216166 114938 216208 115174
rect 215888 114854 216208 114938
rect 215888 114618 215930 114854
rect 216166 114618 216208 114854
rect 215888 114586 216208 114618
rect 207834 100938 207866 101494
rect 208422 100938 208454 101494
rect 207834 65494 208454 100938
rect 217794 111454 218414 146898
rect 217794 110898 217826 111454
rect 218382 110898 218414 111454
rect 215888 79174 216208 79206
rect 215888 78938 215930 79174
rect 216166 78938 216208 79174
rect 215888 78854 216208 78938
rect 215888 78618 215930 78854
rect 216166 78618 216208 78854
rect 215888 78586 216208 78618
rect 207834 64938 207866 65494
rect 208422 64938 208454 65494
rect 207834 29494 208454 64938
rect 217794 75454 218414 110898
rect 217794 74898 217826 75454
rect 218382 74898 218414 75454
rect 215888 43174 216208 43206
rect 215888 42938 215930 43174
rect 216166 42938 216208 43174
rect 215888 42854 216208 42938
rect 215888 42618 215930 42854
rect 216166 42618 216208 42854
rect 215888 42586 216208 42618
rect 207834 28938 207866 29494
rect 208422 28938 208454 29494
rect 207834 -7066 208454 28938
rect 217794 39454 218414 74898
rect 217794 38898 217826 39454
rect 218382 38898 218414 39454
rect 215888 7174 216208 7206
rect 215888 6938 215930 7174
rect 216166 6938 216208 7174
rect 215888 6854 216208 6938
rect 215888 6618 215930 6854
rect 216166 6618 216208 6854
rect 215888 6586 216208 6618
rect 207834 -7622 207866 -7066
rect 208422 -7622 208454 -7066
rect 207834 -7654 208454 -7622
rect 217794 3454 218414 38898
rect 217794 2898 217826 3454
rect 218382 2898 218414 3454
rect 217794 -346 218414 2898
rect 217794 -902 217826 -346
rect 218382 -902 218414 -346
rect 217794 -7654 218414 -902
rect 221514 705798 222134 711590
rect 221514 705242 221546 705798
rect 222102 705242 222134 705798
rect 221514 691174 222134 705242
rect 221514 690618 221546 691174
rect 222102 690618 222134 691174
rect 221514 655174 222134 690618
rect 221514 654618 221546 655174
rect 222102 654618 222134 655174
rect 221514 619174 222134 654618
rect 221514 618618 221546 619174
rect 222102 618618 222134 619174
rect 221514 583174 222134 618618
rect 221514 582618 221546 583174
rect 222102 582618 222134 583174
rect 221514 547174 222134 582618
rect 221514 546618 221546 547174
rect 222102 546618 222134 547174
rect 221514 511174 222134 546618
rect 221514 510618 221546 511174
rect 222102 510618 222134 511174
rect 221514 475174 222134 510618
rect 221514 474618 221546 475174
rect 222102 474618 222134 475174
rect 221514 439174 222134 474618
rect 221514 438618 221546 439174
rect 222102 438618 222134 439174
rect 221514 403174 222134 438618
rect 221514 402618 221546 403174
rect 222102 402618 222134 403174
rect 221514 367174 222134 402618
rect 221514 366618 221546 367174
rect 222102 366618 222134 367174
rect 221514 331174 222134 366618
rect 221514 330618 221546 331174
rect 222102 330618 222134 331174
rect 221514 295174 222134 330618
rect 221514 294618 221546 295174
rect 222102 294618 222134 295174
rect 221514 259174 222134 294618
rect 221514 258618 221546 259174
rect 222102 258618 222134 259174
rect 221514 223174 222134 258618
rect 221514 222618 221546 223174
rect 222102 222618 222134 223174
rect 221514 187174 222134 222618
rect 221514 186618 221546 187174
rect 222102 186618 222134 187174
rect 221514 151174 222134 186618
rect 221514 150618 221546 151174
rect 222102 150618 222134 151174
rect 221514 115174 222134 150618
rect 221514 114618 221546 115174
rect 222102 114618 222134 115174
rect 221514 79174 222134 114618
rect 221514 78618 221546 79174
rect 222102 78618 222134 79174
rect 221514 43174 222134 78618
rect 221514 42618 221546 43174
rect 222102 42618 222134 43174
rect 221514 7174 222134 42618
rect 221514 6618 221546 7174
rect 222102 6618 222134 7174
rect 221514 -1306 222134 6618
rect 221514 -1862 221546 -1306
rect 222102 -1862 222134 -1306
rect 221514 -7654 222134 -1862
rect 225234 706758 225854 711590
rect 225234 706202 225266 706758
rect 225822 706202 225854 706758
rect 225234 694894 225854 706202
rect 225234 694338 225266 694894
rect 225822 694338 225854 694894
rect 225234 658894 225854 694338
rect 225234 658338 225266 658894
rect 225822 658338 225854 658894
rect 225234 622894 225854 658338
rect 225234 622338 225266 622894
rect 225822 622338 225854 622894
rect 225234 586894 225854 622338
rect 225234 586338 225266 586894
rect 225822 586338 225854 586894
rect 225234 550894 225854 586338
rect 225234 550338 225266 550894
rect 225822 550338 225854 550894
rect 225234 514894 225854 550338
rect 225234 514338 225266 514894
rect 225822 514338 225854 514894
rect 225234 478894 225854 514338
rect 225234 478338 225266 478894
rect 225822 478338 225854 478894
rect 225234 442894 225854 478338
rect 225234 442338 225266 442894
rect 225822 442338 225854 442894
rect 225234 406894 225854 442338
rect 225234 406338 225266 406894
rect 225822 406338 225854 406894
rect 225234 370894 225854 406338
rect 225234 370338 225266 370894
rect 225822 370338 225854 370894
rect 225234 334894 225854 370338
rect 225234 334338 225266 334894
rect 225822 334338 225854 334894
rect 225234 298894 225854 334338
rect 225234 298338 225266 298894
rect 225822 298338 225854 298894
rect 225234 262894 225854 298338
rect 225234 262338 225266 262894
rect 225822 262338 225854 262894
rect 225234 226894 225854 262338
rect 225234 226338 225266 226894
rect 225822 226338 225854 226894
rect 225234 190894 225854 226338
rect 225234 190338 225266 190894
rect 225822 190338 225854 190894
rect 225234 154894 225854 190338
rect 225234 154338 225266 154894
rect 225822 154338 225854 154894
rect 225234 118894 225854 154338
rect 225234 118338 225266 118894
rect 225822 118338 225854 118894
rect 225234 82894 225854 118338
rect 225234 82338 225266 82894
rect 225822 82338 225854 82894
rect 225234 46894 225854 82338
rect 225234 46338 225266 46894
rect 225822 46338 225854 46894
rect 225234 10894 225854 46338
rect 225234 10338 225266 10894
rect 225822 10338 225854 10894
rect 225234 -2266 225854 10338
rect 225234 -2822 225266 -2266
rect 225822 -2822 225854 -2266
rect 225234 -7654 225854 -2822
rect 228954 707718 229574 711590
rect 228954 707162 228986 707718
rect 229542 707162 229574 707718
rect 228954 698614 229574 707162
rect 228954 698058 228986 698614
rect 229542 698058 229574 698614
rect 228954 662614 229574 698058
rect 228954 662058 228986 662614
rect 229542 662058 229574 662614
rect 228954 626614 229574 662058
rect 228954 626058 228986 626614
rect 229542 626058 229574 626614
rect 228954 590614 229574 626058
rect 228954 590058 228986 590614
rect 229542 590058 229574 590614
rect 228954 554614 229574 590058
rect 228954 554058 228986 554614
rect 229542 554058 229574 554614
rect 228954 518614 229574 554058
rect 228954 518058 228986 518614
rect 229542 518058 229574 518614
rect 228954 482614 229574 518058
rect 228954 482058 228986 482614
rect 229542 482058 229574 482614
rect 228954 446614 229574 482058
rect 228954 446058 228986 446614
rect 229542 446058 229574 446614
rect 228954 410614 229574 446058
rect 228954 410058 228986 410614
rect 229542 410058 229574 410614
rect 228954 374614 229574 410058
rect 228954 374058 228986 374614
rect 229542 374058 229574 374614
rect 228954 338614 229574 374058
rect 228954 338058 228986 338614
rect 229542 338058 229574 338614
rect 228954 302614 229574 338058
rect 232674 708678 233294 711590
rect 232674 708122 232706 708678
rect 233262 708122 233294 708678
rect 232674 666334 233294 708122
rect 232674 665778 232706 666334
rect 233262 665778 233294 666334
rect 232674 630334 233294 665778
rect 232674 629778 232706 630334
rect 233262 629778 233294 630334
rect 232674 594334 233294 629778
rect 232674 593778 232706 594334
rect 233262 593778 233294 594334
rect 232674 558334 233294 593778
rect 232674 557778 232706 558334
rect 233262 557778 233294 558334
rect 232674 522334 233294 557778
rect 232674 521778 232706 522334
rect 233262 521778 233294 522334
rect 232674 486334 233294 521778
rect 232674 485778 232706 486334
rect 233262 485778 233294 486334
rect 232674 450334 233294 485778
rect 232674 449778 232706 450334
rect 233262 449778 233294 450334
rect 232674 414334 233294 449778
rect 232674 413778 232706 414334
rect 233262 413778 233294 414334
rect 232674 378334 233294 413778
rect 232674 377778 232706 378334
rect 233262 377778 233294 378334
rect 232674 342334 233294 377778
rect 232674 341778 232706 342334
rect 233262 341778 233294 342334
rect 231248 327454 231568 327486
rect 231248 327218 231290 327454
rect 231526 327218 231568 327454
rect 231248 327134 231568 327218
rect 231248 326898 231290 327134
rect 231526 326898 231568 327134
rect 231248 326866 231568 326898
rect 228954 302058 228986 302614
rect 229542 302058 229574 302614
rect 228954 266614 229574 302058
rect 232674 306334 233294 341778
rect 232674 305778 232706 306334
rect 233262 305778 233294 306334
rect 231248 291454 231568 291486
rect 231248 291218 231290 291454
rect 231526 291218 231568 291454
rect 231248 291134 231568 291218
rect 231248 290898 231290 291134
rect 231526 290898 231568 291134
rect 231248 290866 231568 290898
rect 228954 266058 228986 266614
rect 229542 266058 229574 266614
rect 228954 230614 229574 266058
rect 232674 270334 233294 305778
rect 232674 269778 232706 270334
rect 233262 269778 233294 270334
rect 231248 255454 231568 255486
rect 231248 255218 231290 255454
rect 231526 255218 231568 255454
rect 231248 255134 231568 255218
rect 231248 254898 231290 255134
rect 231526 254898 231568 255134
rect 231248 254866 231568 254898
rect 228954 230058 228986 230614
rect 229542 230058 229574 230614
rect 228954 194614 229574 230058
rect 232674 234334 233294 269778
rect 232674 233778 232706 234334
rect 233262 233778 233294 234334
rect 231248 219454 231568 219486
rect 231248 219218 231290 219454
rect 231526 219218 231568 219454
rect 231248 219134 231568 219218
rect 231248 218898 231290 219134
rect 231526 218898 231568 219134
rect 231248 218866 231568 218898
rect 228954 194058 228986 194614
rect 229542 194058 229574 194614
rect 228954 158614 229574 194058
rect 232674 198334 233294 233778
rect 232674 197778 232706 198334
rect 233262 197778 233294 198334
rect 231248 183454 231568 183486
rect 231248 183218 231290 183454
rect 231526 183218 231568 183454
rect 231248 183134 231568 183218
rect 231248 182898 231290 183134
rect 231526 182898 231568 183134
rect 231248 182866 231568 182898
rect 228954 158058 228986 158614
rect 229542 158058 229574 158614
rect 228954 122614 229574 158058
rect 232674 162334 233294 197778
rect 232674 161778 232706 162334
rect 233262 161778 233294 162334
rect 231248 147454 231568 147486
rect 231248 147218 231290 147454
rect 231526 147218 231568 147454
rect 231248 147134 231568 147218
rect 231248 146898 231290 147134
rect 231526 146898 231568 147134
rect 231248 146866 231568 146898
rect 228954 122058 228986 122614
rect 229542 122058 229574 122614
rect 228954 86614 229574 122058
rect 232674 126334 233294 161778
rect 232674 125778 232706 126334
rect 233262 125778 233294 126334
rect 231248 111454 231568 111486
rect 231248 111218 231290 111454
rect 231526 111218 231568 111454
rect 231248 111134 231568 111218
rect 231248 110898 231290 111134
rect 231526 110898 231568 111134
rect 231248 110866 231568 110898
rect 228954 86058 228986 86614
rect 229542 86058 229574 86614
rect 228954 50614 229574 86058
rect 232674 90334 233294 125778
rect 232674 89778 232706 90334
rect 233262 89778 233294 90334
rect 231248 75454 231568 75486
rect 231248 75218 231290 75454
rect 231526 75218 231568 75454
rect 231248 75134 231568 75218
rect 231248 74898 231290 75134
rect 231526 74898 231568 75134
rect 231248 74866 231568 74898
rect 228954 50058 228986 50614
rect 229542 50058 229574 50614
rect 228954 14614 229574 50058
rect 232674 54334 233294 89778
rect 232674 53778 232706 54334
rect 233262 53778 233294 54334
rect 231248 39454 231568 39486
rect 231248 39218 231290 39454
rect 231526 39218 231568 39454
rect 231248 39134 231568 39218
rect 231248 38898 231290 39134
rect 231526 38898 231568 39134
rect 231248 38866 231568 38898
rect 228954 14058 228986 14614
rect 229542 14058 229574 14614
rect 228954 -3226 229574 14058
rect 228954 -3782 228986 -3226
rect 229542 -3782 229574 -3226
rect 228954 -7654 229574 -3782
rect 232674 18334 233294 53778
rect 232674 17778 232706 18334
rect 233262 17778 233294 18334
rect 232674 -4186 233294 17778
rect 232674 -4742 232706 -4186
rect 233262 -4742 233294 -4186
rect 232674 -7654 233294 -4742
rect 236394 709638 237014 711590
rect 236394 709082 236426 709638
rect 236982 709082 237014 709638
rect 236394 670054 237014 709082
rect 236394 669498 236426 670054
rect 236982 669498 237014 670054
rect 236394 634054 237014 669498
rect 236394 633498 236426 634054
rect 236982 633498 237014 634054
rect 236394 598054 237014 633498
rect 236394 597498 236426 598054
rect 236982 597498 237014 598054
rect 236394 562054 237014 597498
rect 236394 561498 236426 562054
rect 236982 561498 237014 562054
rect 236394 526054 237014 561498
rect 236394 525498 236426 526054
rect 236982 525498 237014 526054
rect 236394 490054 237014 525498
rect 236394 489498 236426 490054
rect 236982 489498 237014 490054
rect 236394 454054 237014 489498
rect 236394 453498 236426 454054
rect 236982 453498 237014 454054
rect 236394 418054 237014 453498
rect 236394 417498 236426 418054
rect 236982 417498 237014 418054
rect 236394 382054 237014 417498
rect 236394 381498 236426 382054
rect 236982 381498 237014 382054
rect 236394 346054 237014 381498
rect 236394 345498 236426 346054
rect 236982 345498 237014 346054
rect 236394 310054 237014 345498
rect 236394 309498 236426 310054
rect 236982 309498 237014 310054
rect 236394 274054 237014 309498
rect 236394 273498 236426 274054
rect 236982 273498 237014 274054
rect 236394 238054 237014 273498
rect 236394 237498 236426 238054
rect 236982 237498 237014 238054
rect 236394 202054 237014 237498
rect 236394 201498 236426 202054
rect 236982 201498 237014 202054
rect 236394 166054 237014 201498
rect 236394 165498 236426 166054
rect 236982 165498 237014 166054
rect 236394 130054 237014 165498
rect 236394 129498 236426 130054
rect 236982 129498 237014 130054
rect 236394 94054 237014 129498
rect 236394 93498 236426 94054
rect 236982 93498 237014 94054
rect 236394 58054 237014 93498
rect 236394 57498 236426 58054
rect 236982 57498 237014 58054
rect 236394 22054 237014 57498
rect 240114 710598 240734 711590
rect 240114 710042 240146 710598
rect 240702 710042 240734 710598
rect 240114 673774 240734 710042
rect 240114 673218 240146 673774
rect 240702 673218 240734 673774
rect 240114 637774 240734 673218
rect 240114 637218 240146 637774
rect 240702 637218 240734 637774
rect 240114 601774 240734 637218
rect 240114 601218 240146 601774
rect 240702 601218 240734 601774
rect 240114 565774 240734 601218
rect 240114 565218 240146 565774
rect 240702 565218 240734 565774
rect 240114 529774 240734 565218
rect 240114 529218 240146 529774
rect 240702 529218 240734 529774
rect 240114 493774 240734 529218
rect 240114 493218 240146 493774
rect 240702 493218 240734 493774
rect 240114 457774 240734 493218
rect 240114 457218 240146 457774
rect 240702 457218 240734 457774
rect 240114 421774 240734 457218
rect 240114 421218 240146 421774
rect 240702 421218 240734 421774
rect 240114 385774 240734 421218
rect 240114 385218 240146 385774
rect 240702 385218 240734 385774
rect 240114 349774 240734 385218
rect 240114 349218 240146 349774
rect 240702 349218 240734 349774
rect 240114 313774 240734 349218
rect 240114 313218 240146 313774
rect 240702 313218 240734 313774
rect 240114 277774 240734 313218
rect 240114 277218 240146 277774
rect 240702 277218 240734 277774
rect 240114 241774 240734 277218
rect 240114 241218 240146 241774
rect 240702 241218 240734 241774
rect 240114 205774 240734 241218
rect 240114 205218 240146 205774
rect 240702 205218 240734 205774
rect 240114 169774 240734 205218
rect 240114 169218 240146 169774
rect 240702 169218 240734 169774
rect 240114 133774 240734 169218
rect 240114 133218 240146 133774
rect 240702 133218 240734 133774
rect 240114 97774 240734 133218
rect 240114 97218 240146 97774
rect 240702 97218 240734 97774
rect 240114 61774 240734 97218
rect 240114 61218 240146 61774
rect 240702 61218 240734 61774
rect 240114 27193 240734 61218
rect 243834 711558 244454 711590
rect 243834 711002 243866 711558
rect 244422 711002 244454 711558
rect 243834 677494 244454 711002
rect 243834 676938 243866 677494
rect 244422 676938 244454 677494
rect 243834 641494 244454 676938
rect 243834 640938 243866 641494
rect 244422 640938 244454 641494
rect 243834 605494 244454 640938
rect 243834 604938 243866 605494
rect 244422 604938 244454 605494
rect 243834 569494 244454 604938
rect 243834 568938 243866 569494
rect 244422 568938 244454 569494
rect 243834 533494 244454 568938
rect 243834 532938 243866 533494
rect 244422 532938 244454 533494
rect 243834 497494 244454 532938
rect 243834 496938 243866 497494
rect 244422 496938 244454 497494
rect 243834 461494 244454 496938
rect 243834 460938 243866 461494
rect 244422 460938 244454 461494
rect 243834 425494 244454 460938
rect 243834 424938 243866 425494
rect 244422 424938 244454 425494
rect 243834 389494 244454 424938
rect 243834 388938 243866 389494
rect 244422 388938 244454 389494
rect 243834 353494 244454 388938
rect 243834 352938 243866 353494
rect 244422 352938 244454 353494
rect 243834 317494 244454 352938
rect 253794 704838 254414 711590
rect 253794 704282 253826 704838
rect 254382 704282 254414 704838
rect 253794 687454 254414 704282
rect 253794 686898 253826 687454
rect 254382 686898 254414 687454
rect 253794 651454 254414 686898
rect 253794 650898 253826 651454
rect 254382 650898 254414 651454
rect 253794 615454 254414 650898
rect 253794 614898 253826 615454
rect 254382 614898 254414 615454
rect 253794 579454 254414 614898
rect 253794 578898 253826 579454
rect 254382 578898 254414 579454
rect 253794 543454 254414 578898
rect 253794 542898 253826 543454
rect 254382 542898 254414 543454
rect 253794 507454 254414 542898
rect 253794 506898 253826 507454
rect 254382 506898 254414 507454
rect 253794 471454 254414 506898
rect 253794 470898 253826 471454
rect 254382 470898 254414 471454
rect 253794 435454 254414 470898
rect 253794 434898 253826 435454
rect 254382 434898 254414 435454
rect 253794 399454 254414 434898
rect 253794 398898 253826 399454
rect 254382 398898 254414 399454
rect 253794 363454 254414 398898
rect 253794 362898 253826 363454
rect 254382 362898 254414 363454
rect 246608 331174 246928 331206
rect 246608 330938 246650 331174
rect 246886 330938 246928 331174
rect 246608 330854 246928 330938
rect 246608 330618 246650 330854
rect 246886 330618 246928 330854
rect 246608 330586 246928 330618
rect 243834 316938 243866 317494
rect 244422 316938 244454 317494
rect 243834 281494 244454 316938
rect 253794 327454 254414 362898
rect 253794 326898 253826 327454
rect 254382 326898 254414 327454
rect 246608 295174 246928 295206
rect 246608 294938 246650 295174
rect 246886 294938 246928 295174
rect 246608 294854 246928 294938
rect 246608 294618 246650 294854
rect 246886 294618 246928 294854
rect 246608 294586 246928 294618
rect 243834 280938 243866 281494
rect 244422 280938 244454 281494
rect 243834 245494 244454 280938
rect 253794 291454 254414 326898
rect 253794 290898 253826 291454
rect 254382 290898 254414 291454
rect 246608 259174 246928 259206
rect 246608 258938 246650 259174
rect 246886 258938 246928 259174
rect 246608 258854 246928 258938
rect 246608 258618 246650 258854
rect 246886 258618 246928 258854
rect 246608 258586 246928 258618
rect 243834 244938 243866 245494
rect 244422 244938 244454 245494
rect 243834 209494 244454 244938
rect 253794 255454 254414 290898
rect 253794 254898 253826 255454
rect 254382 254898 254414 255454
rect 246608 223174 246928 223206
rect 246608 222938 246650 223174
rect 246886 222938 246928 223174
rect 246608 222854 246928 222938
rect 246608 222618 246650 222854
rect 246886 222618 246928 222854
rect 246608 222586 246928 222618
rect 243834 208938 243866 209494
rect 244422 208938 244454 209494
rect 243834 173494 244454 208938
rect 253794 219454 254414 254898
rect 253794 218898 253826 219454
rect 254382 218898 254414 219454
rect 246608 187174 246928 187206
rect 246608 186938 246650 187174
rect 246886 186938 246928 187174
rect 246608 186854 246928 186938
rect 246608 186618 246650 186854
rect 246886 186618 246928 186854
rect 246608 186586 246928 186618
rect 243834 172938 243866 173494
rect 244422 172938 244454 173494
rect 243834 137494 244454 172938
rect 253794 183454 254414 218898
rect 253794 182898 253826 183454
rect 254382 182898 254414 183454
rect 246608 151174 246928 151206
rect 246608 150938 246650 151174
rect 246886 150938 246928 151174
rect 246608 150854 246928 150938
rect 246608 150618 246650 150854
rect 246886 150618 246928 150854
rect 246608 150586 246928 150618
rect 243834 136938 243866 137494
rect 244422 136938 244454 137494
rect 243834 101494 244454 136938
rect 253794 147454 254414 182898
rect 253794 146898 253826 147454
rect 254382 146898 254414 147454
rect 246608 115174 246928 115206
rect 246608 114938 246650 115174
rect 246886 114938 246928 115174
rect 246608 114854 246928 114938
rect 246608 114618 246650 114854
rect 246886 114618 246928 114854
rect 246608 114586 246928 114618
rect 243834 100938 243866 101494
rect 244422 100938 244454 101494
rect 243834 65494 244454 100938
rect 253794 111454 254414 146898
rect 253794 110898 253826 111454
rect 254382 110898 254414 111454
rect 246608 79174 246928 79206
rect 246608 78938 246650 79174
rect 246886 78938 246928 79174
rect 246608 78854 246928 78938
rect 246608 78618 246650 78854
rect 246886 78618 246928 78854
rect 246608 78586 246928 78618
rect 243834 64938 243866 65494
rect 244422 64938 244454 65494
rect 243834 29494 244454 64938
rect 253794 75454 254414 110898
rect 253794 74898 253826 75454
rect 254382 74898 254414 75454
rect 246608 43174 246928 43206
rect 246608 42938 246650 43174
rect 246886 42938 246928 43174
rect 246608 42854 246928 42938
rect 246608 42618 246650 42854
rect 246886 42618 246928 42854
rect 246608 42586 246928 42618
rect 243834 28938 243866 29494
rect 244422 28938 244454 29494
rect 243834 27193 244454 28938
rect 253794 39454 254414 74898
rect 253794 38898 253826 39454
rect 254382 38898 254414 39454
rect 253794 27193 254414 38898
rect 257514 705798 258134 711590
rect 257514 705242 257546 705798
rect 258102 705242 258134 705798
rect 257514 691174 258134 705242
rect 257514 690618 257546 691174
rect 258102 690618 258134 691174
rect 257514 655174 258134 690618
rect 257514 654618 257546 655174
rect 258102 654618 258134 655174
rect 257514 619174 258134 654618
rect 257514 618618 257546 619174
rect 258102 618618 258134 619174
rect 257514 583174 258134 618618
rect 257514 582618 257546 583174
rect 258102 582618 258134 583174
rect 257514 547174 258134 582618
rect 257514 546618 257546 547174
rect 258102 546618 258134 547174
rect 257514 511174 258134 546618
rect 257514 510618 257546 511174
rect 258102 510618 258134 511174
rect 257514 475174 258134 510618
rect 257514 474618 257546 475174
rect 258102 474618 258134 475174
rect 257514 439174 258134 474618
rect 257514 438618 257546 439174
rect 258102 438618 258134 439174
rect 257514 403174 258134 438618
rect 257514 402618 257546 403174
rect 258102 402618 258134 403174
rect 257514 367174 258134 402618
rect 257514 366618 257546 367174
rect 258102 366618 258134 367174
rect 257514 331174 258134 366618
rect 257514 330618 257546 331174
rect 258102 330618 258134 331174
rect 257514 295174 258134 330618
rect 257514 294618 257546 295174
rect 258102 294618 258134 295174
rect 257514 259174 258134 294618
rect 257514 258618 257546 259174
rect 258102 258618 258134 259174
rect 257514 223174 258134 258618
rect 257514 222618 257546 223174
rect 258102 222618 258134 223174
rect 257514 187174 258134 222618
rect 257514 186618 257546 187174
rect 258102 186618 258134 187174
rect 257514 151174 258134 186618
rect 257514 150618 257546 151174
rect 258102 150618 258134 151174
rect 257514 115174 258134 150618
rect 257514 114618 257546 115174
rect 258102 114618 258134 115174
rect 257514 79174 258134 114618
rect 257514 78618 257546 79174
rect 258102 78618 258134 79174
rect 257514 43174 258134 78618
rect 257514 42618 257546 43174
rect 258102 42618 258134 43174
rect 257514 27193 258134 42618
rect 261234 706758 261854 711590
rect 261234 706202 261266 706758
rect 261822 706202 261854 706758
rect 261234 694894 261854 706202
rect 261234 694338 261266 694894
rect 261822 694338 261854 694894
rect 261234 658894 261854 694338
rect 261234 658338 261266 658894
rect 261822 658338 261854 658894
rect 261234 622894 261854 658338
rect 261234 622338 261266 622894
rect 261822 622338 261854 622894
rect 261234 586894 261854 622338
rect 261234 586338 261266 586894
rect 261822 586338 261854 586894
rect 261234 550894 261854 586338
rect 261234 550338 261266 550894
rect 261822 550338 261854 550894
rect 261234 514894 261854 550338
rect 261234 514338 261266 514894
rect 261822 514338 261854 514894
rect 261234 478894 261854 514338
rect 261234 478338 261266 478894
rect 261822 478338 261854 478894
rect 261234 442894 261854 478338
rect 261234 442338 261266 442894
rect 261822 442338 261854 442894
rect 261234 406894 261854 442338
rect 261234 406338 261266 406894
rect 261822 406338 261854 406894
rect 261234 370894 261854 406338
rect 261234 370338 261266 370894
rect 261822 370338 261854 370894
rect 261234 334894 261854 370338
rect 261234 334338 261266 334894
rect 261822 334338 261854 334894
rect 261234 298894 261854 334338
rect 264954 707718 265574 711590
rect 264954 707162 264986 707718
rect 265542 707162 265574 707718
rect 264954 698614 265574 707162
rect 264954 698058 264986 698614
rect 265542 698058 265574 698614
rect 264954 662614 265574 698058
rect 264954 662058 264986 662614
rect 265542 662058 265574 662614
rect 264954 626614 265574 662058
rect 264954 626058 264986 626614
rect 265542 626058 265574 626614
rect 264954 590614 265574 626058
rect 264954 590058 264986 590614
rect 265542 590058 265574 590614
rect 264954 554614 265574 590058
rect 264954 554058 264986 554614
rect 265542 554058 265574 554614
rect 264954 518614 265574 554058
rect 264954 518058 264986 518614
rect 265542 518058 265574 518614
rect 264954 482614 265574 518058
rect 264954 482058 264986 482614
rect 265542 482058 265574 482614
rect 264954 446614 265574 482058
rect 264954 446058 264986 446614
rect 265542 446058 265574 446614
rect 264954 410614 265574 446058
rect 264954 410058 264986 410614
rect 265542 410058 265574 410614
rect 264954 374614 265574 410058
rect 264954 374058 264986 374614
rect 265542 374058 265574 374614
rect 264954 338614 265574 374058
rect 264954 338058 264986 338614
rect 265542 338058 265574 338614
rect 261968 327454 262288 327486
rect 261968 327218 262010 327454
rect 262246 327218 262288 327454
rect 261968 327134 262288 327218
rect 261968 326898 262010 327134
rect 262246 326898 262288 327134
rect 261968 326866 262288 326898
rect 261234 298338 261266 298894
rect 261822 298338 261854 298894
rect 261234 262894 261854 298338
rect 264954 302614 265574 338058
rect 264954 302058 264986 302614
rect 265542 302058 265574 302614
rect 261968 291454 262288 291486
rect 261968 291218 262010 291454
rect 262246 291218 262288 291454
rect 261968 291134 262288 291218
rect 261968 290898 262010 291134
rect 262246 290898 262288 291134
rect 261968 290866 262288 290898
rect 261234 262338 261266 262894
rect 261822 262338 261854 262894
rect 261234 226894 261854 262338
rect 264954 266614 265574 302058
rect 264954 266058 264986 266614
rect 265542 266058 265574 266614
rect 261968 255454 262288 255486
rect 261968 255218 262010 255454
rect 262246 255218 262288 255454
rect 261968 255134 262288 255218
rect 261968 254898 262010 255134
rect 262246 254898 262288 255134
rect 261968 254866 262288 254898
rect 261234 226338 261266 226894
rect 261822 226338 261854 226894
rect 261234 190894 261854 226338
rect 264954 230614 265574 266058
rect 264954 230058 264986 230614
rect 265542 230058 265574 230614
rect 261968 219454 262288 219486
rect 261968 219218 262010 219454
rect 262246 219218 262288 219454
rect 261968 219134 262288 219218
rect 261968 218898 262010 219134
rect 262246 218898 262288 219134
rect 261968 218866 262288 218898
rect 261234 190338 261266 190894
rect 261822 190338 261854 190894
rect 261234 154894 261854 190338
rect 264954 194614 265574 230058
rect 264954 194058 264986 194614
rect 265542 194058 265574 194614
rect 261968 183454 262288 183486
rect 261968 183218 262010 183454
rect 262246 183218 262288 183454
rect 261968 183134 262288 183218
rect 261968 182898 262010 183134
rect 262246 182898 262288 183134
rect 261968 182866 262288 182898
rect 261234 154338 261266 154894
rect 261822 154338 261854 154894
rect 261234 118894 261854 154338
rect 264954 158614 265574 194058
rect 264954 158058 264986 158614
rect 265542 158058 265574 158614
rect 261968 147454 262288 147486
rect 261968 147218 262010 147454
rect 262246 147218 262288 147454
rect 261968 147134 262288 147218
rect 261968 146898 262010 147134
rect 262246 146898 262288 147134
rect 261968 146866 262288 146898
rect 261234 118338 261266 118894
rect 261822 118338 261854 118894
rect 261234 82894 261854 118338
rect 264954 122614 265574 158058
rect 264954 122058 264986 122614
rect 265542 122058 265574 122614
rect 261968 111454 262288 111486
rect 261968 111218 262010 111454
rect 262246 111218 262288 111454
rect 261968 111134 262288 111218
rect 261968 110898 262010 111134
rect 262246 110898 262288 111134
rect 261968 110866 262288 110898
rect 261234 82338 261266 82894
rect 261822 82338 261854 82894
rect 261234 46894 261854 82338
rect 264954 86614 265574 122058
rect 264954 86058 264986 86614
rect 265542 86058 265574 86614
rect 261968 75454 262288 75486
rect 261968 75218 262010 75454
rect 262246 75218 262288 75454
rect 261968 75134 262288 75218
rect 261968 74898 262010 75134
rect 262246 74898 262288 75134
rect 261968 74866 262288 74898
rect 261234 46338 261266 46894
rect 261822 46338 261854 46894
rect 236394 21498 236426 22054
rect 236982 21498 237014 22054
rect 236394 -5146 237014 21498
rect 261234 10894 261854 46338
rect 264954 50614 265574 86058
rect 264954 50058 264986 50614
rect 265542 50058 265574 50614
rect 261968 39454 262288 39486
rect 261968 39218 262010 39454
rect 262246 39218 262288 39454
rect 261968 39134 262288 39218
rect 261968 38898 262010 39134
rect 262246 38898 262288 39134
rect 261968 38866 262288 38898
rect 261234 10338 261266 10894
rect 261822 10338 261854 10894
rect 246608 7174 246928 7206
rect 246608 6938 246650 7174
rect 246886 6938 246928 7174
rect 246608 6854 246928 6938
rect 246608 6618 246650 6854
rect 246886 6618 246928 6854
rect 246608 6586 246928 6618
rect 236394 -5702 236426 -5146
rect 236982 -5702 237014 -5146
rect 236394 -7654 237014 -5702
rect 253794 3454 254414 4103
rect 253794 2898 253826 3454
rect 254382 2898 254414 3454
rect 253794 -346 254414 2898
rect 253794 -902 253826 -346
rect 254382 -902 254414 -346
rect 253794 -7654 254414 -902
rect 261234 -2266 261854 10338
rect 261234 -2822 261266 -2266
rect 261822 -2822 261854 -2266
rect 261234 -7654 261854 -2822
rect 264954 14614 265574 50058
rect 264954 14058 264986 14614
rect 265542 14058 265574 14614
rect 264954 -3226 265574 14058
rect 264954 -3782 264986 -3226
rect 265542 -3782 265574 -3226
rect 264954 -7654 265574 -3782
rect 268674 708678 269294 711590
rect 268674 708122 268706 708678
rect 269262 708122 269294 708678
rect 268674 666334 269294 708122
rect 268674 665778 268706 666334
rect 269262 665778 269294 666334
rect 268674 630334 269294 665778
rect 268674 629778 268706 630334
rect 269262 629778 269294 630334
rect 268674 594334 269294 629778
rect 268674 593778 268706 594334
rect 269262 593778 269294 594334
rect 268674 558334 269294 593778
rect 268674 557778 268706 558334
rect 269262 557778 269294 558334
rect 268674 522334 269294 557778
rect 268674 521778 268706 522334
rect 269262 521778 269294 522334
rect 268674 486334 269294 521778
rect 268674 485778 268706 486334
rect 269262 485778 269294 486334
rect 268674 450334 269294 485778
rect 268674 449778 268706 450334
rect 269262 449778 269294 450334
rect 268674 414334 269294 449778
rect 268674 413778 268706 414334
rect 269262 413778 269294 414334
rect 268674 378334 269294 413778
rect 268674 377778 268706 378334
rect 269262 377778 269294 378334
rect 268674 342334 269294 377778
rect 268674 341778 268706 342334
rect 269262 341778 269294 342334
rect 268674 306334 269294 341778
rect 268674 305778 268706 306334
rect 269262 305778 269294 306334
rect 268674 270334 269294 305778
rect 268674 269778 268706 270334
rect 269262 269778 269294 270334
rect 268674 234334 269294 269778
rect 268674 233778 268706 234334
rect 269262 233778 269294 234334
rect 268674 198334 269294 233778
rect 268674 197778 268706 198334
rect 269262 197778 269294 198334
rect 268674 162334 269294 197778
rect 268674 161778 268706 162334
rect 269262 161778 269294 162334
rect 268674 126334 269294 161778
rect 268674 125778 268706 126334
rect 269262 125778 269294 126334
rect 268674 90334 269294 125778
rect 268674 89778 268706 90334
rect 269262 89778 269294 90334
rect 268674 54334 269294 89778
rect 268674 53778 268706 54334
rect 269262 53778 269294 54334
rect 268674 18334 269294 53778
rect 268674 17778 268706 18334
rect 269262 17778 269294 18334
rect 268674 -4186 269294 17778
rect 268674 -4742 268706 -4186
rect 269262 -4742 269294 -4186
rect 268674 -7654 269294 -4742
rect 272394 709638 273014 711590
rect 272394 709082 272426 709638
rect 272982 709082 273014 709638
rect 272394 670054 273014 709082
rect 272394 669498 272426 670054
rect 272982 669498 273014 670054
rect 272394 634054 273014 669498
rect 272394 633498 272426 634054
rect 272982 633498 273014 634054
rect 272394 598054 273014 633498
rect 272394 597498 272426 598054
rect 272982 597498 273014 598054
rect 272394 562054 273014 597498
rect 272394 561498 272426 562054
rect 272982 561498 273014 562054
rect 272394 526054 273014 561498
rect 272394 525498 272426 526054
rect 272982 525498 273014 526054
rect 272394 490054 273014 525498
rect 272394 489498 272426 490054
rect 272982 489498 273014 490054
rect 272394 454054 273014 489498
rect 272394 453498 272426 454054
rect 272982 453498 273014 454054
rect 272394 418054 273014 453498
rect 272394 417498 272426 418054
rect 272982 417498 273014 418054
rect 272394 382054 273014 417498
rect 272394 381498 272426 382054
rect 272982 381498 273014 382054
rect 272394 346054 273014 381498
rect 272394 345498 272426 346054
rect 272982 345498 273014 346054
rect 272394 310054 273014 345498
rect 272394 309498 272426 310054
rect 272982 309498 273014 310054
rect 272394 274054 273014 309498
rect 272394 273498 272426 274054
rect 272982 273498 273014 274054
rect 272394 238054 273014 273498
rect 272394 237498 272426 238054
rect 272982 237498 273014 238054
rect 272394 202054 273014 237498
rect 272394 201498 272426 202054
rect 272982 201498 273014 202054
rect 272394 166054 273014 201498
rect 272394 165498 272426 166054
rect 272982 165498 273014 166054
rect 272394 130054 273014 165498
rect 272394 129498 272426 130054
rect 272982 129498 273014 130054
rect 272394 94054 273014 129498
rect 272394 93498 272426 94054
rect 272982 93498 273014 94054
rect 272394 58054 273014 93498
rect 272394 57498 272426 58054
rect 272982 57498 273014 58054
rect 272394 22054 273014 57498
rect 272394 21498 272426 22054
rect 272982 21498 273014 22054
rect 272394 -5146 273014 21498
rect 272394 -5702 272426 -5146
rect 272982 -5702 273014 -5146
rect 272394 -7654 273014 -5702
rect 276114 710598 276734 711590
rect 276114 710042 276146 710598
rect 276702 710042 276734 710598
rect 276114 673774 276734 710042
rect 276114 673218 276146 673774
rect 276702 673218 276734 673774
rect 276114 637774 276734 673218
rect 276114 637218 276146 637774
rect 276702 637218 276734 637774
rect 276114 601774 276734 637218
rect 276114 601218 276146 601774
rect 276702 601218 276734 601774
rect 276114 565774 276734 601218
rect 276114 565218 276146 565774
rect 276702 565218 276734 565774
rect 276114 529774 276734 565218
rect 276114 529218 276146 529774
rect 276702 529218 276734 529774
rect 276114 493774 276734 529218
rect 276114 493218 276146 493774
rect 276702 493218 276734 493774
rect 276114 457774 276734 493218
rect 276114 457218 276146 457774
rect 276702 457218 276734 457774
rect 276114 421774 276734 457218
rect 276114 421218 276146 421774
rect 276702 421218 276734 421774
rect 276114 385774 276734 421218
rect 276114 385218 276146 385774
rect 276702 385218 276734 385774
rect 276114 349774 276734 385218
rect 276114 349218 276146 349774
rect 276702 349218 276734 349774
rect 276114 313774 276734 349218
rect 279834 711558 280454 711590
rect 279834 711002 279866 711558
rect 280422 711002 280454 711558
rect 279834 677494 280454 711002
rect 279834 676938 279866 677494
rect 280422 676938 280454 677494
rect 279834 641494 280454 676938
rect 279834 640938 279866 641494
rect 280422 640938 280454 641494
rect 279834 605494 280454 640938
rect 279834 604938 279866 605494
rect 280422 604938 280454 605494
rect 279834 569494 280454 604938
rect 279834 568938 279866 569494
rect 280422 568938 280454 569494
rect 279834 533494 280454 568938
rect 279834 532938 279866 533494
rect 280422 532938 280454 533494
rect 279834 497494 280454 532938
rect 279834 496938 279866 497494
rect 280422 496938 280454 497494
rect 279834 461494 280454 496938
rect 279834 460938 279866 461494
rect 280422 460938 280454 461494
rect 279834 425494 280454 460938
rect 279834 424938 279866 425494
rect 280422 424938 280454 425494
rect 279834 389494 280454 424938
rect 279834 388938 279866 389494
rect 280422 388938 280454 389494
rect 279834 353494 280454 388938
rect 279834 352938 279866 353494
rect 280422 352938 280454 353494
rect 277328 331174 277648 331206
rect 277328 330938 277370 331174
rect 277606 330938 277648 331174
rect 277328 330854 277648 330938
rect 277328 330618 277370 330854
rect 277606 330618 277648 330854
rect 277328 330586 277648 330618
rect 276114 313218 276146 313774
rect 276702 313218 276734 313774
rect 276114 277774 276734 313218
rect 279834 317494 280454 352938
rect 279834 316938 279866 317494
rect 280422 316938 280454 317494
rect 277328 295174 277648 295206
rect 277328 294938 277370 295174
rect 277606 294938 277648 295174
rect 277328 294854 277648 294938
rect 277328 294618 277370 294854
rect 277606 294618 277648 294854
rect 277328 294586 277648 294618
rect 276114 277218 276146 277774
rect 276702 277218 276734 277774
rect 276114 241774 276734 277218
rect 279834 281494 280454 316938
rect 279834 280938 279866 281494
rect 280422 280938 280454 281494
rect 277328 259174 277648 259206
rect 277328 258938 277370 259174
rect 277606 258938 277648 259174
rect 277328 258854 277648 258938
rect 277328 258618 277370 258854
rect 277606 258618 277648 258854
rect 277328 258586 277648 258618
rect 276114 241218 276146 241774
rect 276702 241218 276734 241774
rect 276114 205774 276734 241218
rect 279834 245494 280454 280938
rect 279834 244938 279866 245494
rect 280422 244938 280454 245494
rect 277328 223174 277648 223206
rect 277328 222938 277370 223174
rect 277606 222938 277648 223174
rect 277328 222854 277648 222938
rect 277328 222618 277370 222854
rect 277606 222618 277648 222854
rect 277328 222586 277648 222618
rect 276114 205218 276146 205774
rect 276702 205218 276734 205774
rect 276114 169774 276734 205218
rect 279834 209494 280454 244938
rect 279834 208938 279866 209494
rect 280422 208938 280454 209494
rect 277328 187174 277648 187206
rect 277328 186938 277370 187174
rect 277606 186938 277648 187174
rect 277328 186854 277648 186938
rect 277328 186618 277370 186854
rect 277606 186618 277648 186854
rect 277328 186586 277648 186618
rect 276114 169218 276146 169774
rect 276702 169218 276734 169774
rect 276114 133774 276734 169218
rect 279834 173494 280454 208938
rect 279834 172938 279866 173494
rect 280422 172938 280454 173494
rect 277328 151174 277648 151206
rect 277328 150938 277370 151174
rect 277606 150938 277648 151174
rect 277328 150854 277648 150938
rect 277328 150618 277370 150854
rect 277606 150618 277648 150854
rect 277328 150586 277648 150618
rect 276114 133218 276146 133774
rect 276702 133218 276734 133774
rect 276114 97774 276734 133218
rect 279834 137494 280454 172938
rect 279834 136938 279866 137494
rect 280422 136938 280454 137494
rect 277328 115174 277648 115206
rect 277328 114938 277370 115174
rect 277606 114938 277648 115174
rect 277328 114854 277648 114938
rect 277328 114618 277370 114854
rect 277606 114618 277648 114854
rect 277328 114586 277648 114618
rect 276114 97218 276146 97774
rect 276702 97218 276734 97774
rect 276114 61774 276734 97218
rect 279834 101494 280454 136938
rect 279834 100938 279866 101494
rect 280422 100938 280454 101494
rect 277328 79174 277648 79206
rect 277328 78938 277370 79174
rect 277606 78938 277648 79174
rect 277328 78854 277648 78938
rect 277328 78618 277370 78854
rect 277606 78618 277648 78854
rect 277328 78586 277648 78618
rect 276114 61218 276146 61774
rect 276702 61218 276734 61774
rect 276114 25774 276734 61218
rect 279834 65494 280454 100938
rect 279834 64938 279866 65494
rect 280422 64938 280454 65494
rect 277328 43174 277648 43206
rect 277328 42938 277370 43174
rect 277606 42938 277648 43174
rect 277328 42854 277648 42938
rect 277328 42618 277370 42854
rect 277606 42618 277648 42854
rect 277328 42586 277648 42618
rect 276114 25218 276146 25774
rect 276702 25218 276734 25774
rect 276114 -6106 276734 25218
rect 279834 29494 280454 64938
rect 279834 28938 279866 29494
rect 280422 28938 280454 29494
rect 277328 7174 277648 7206
rect 277328 6938 277370 7174
rect 277606 6938 277648 7174
rect 277328 6854 277648 6938
rect 277328 6618 277370 6854
rect 277606 6618 277648 6854
rect 277328 6586 277648 6618
rect 276114 -6662 276146 -6106
rect 276702 -6662 276734 -6106
rect 276114 -7654 276734 -6662
rect 279834 -7066 280454 28938
rect 279834 -7622 279866 -7066
rect 280422 -7622 280454 -7066
rect 279834 -7654 280454 -7622
rect 289794 704838 290414 711590
rect 289794 704282 289826 704838
rect 290382 704282 290414 704838
rect 289794 687454 290414 704282
rect 289794 686898 289826 687454
rect 290382 686898 290414 687454
rect 289794 651454 290414 686898
rect 289794 650898 289826 651454
rect 290382 650898 290414 651454
rect 289794 615454 290414 650898
rect 289794 614898 289826 615454
rect 290382 614898 290414 615454
rect 289794 579454 290414 614898
rect 289794 578898 289826 579454
rect 290382 578898 290414 579454
rect 289794 543454 290414 578898
rect 289794 542898 289826 543454
rect 290382 542898 290414 543454
rect 289794 507454 290414 542898
rect 289794 506898 289826 507454
rect 290382 506898 290414 507454
rect 289794 471454 290414 506898
rect 289794 470898 289826 471454
rect 290382 470898 290414 471454
rect 289794 435454 290414 470898
rect 289794 434898 289826 435454
rect 290382 434898 290414 435454
rect 289794 399454 290414 434898
rect 289794 398898 289826 399454
rect 290382 398898 290414 399454
rect 289794 363454 290414 398898
rect 289794 362898 289826 363454
rect 290382 362898 290414 363454
rect 289794 327454 290414 362898
rect 293514 705798 294134 711590
rect 293514 705242 293546 705798
rect 294102 705242 294134 705798
rect 293514 691174 294134 705242
rect 293514 690618 293546 691174
rect 294102 690618 294134 691174
rect 293514 655174 294134 690618
rect 293514 654618 293546 655174
rect 294102 654618 294134 655174
rect 293514 619174 294134 654618
rect 293514 618618 293546 619174
rect 294102 618618 294134 619174
rect 293514 583174 294134 618618
rect 293514 582618 293546 583174
rect 294102 582618 294134 583174
rect 293514 547174 294134 582618
rect 293514 546618 293546 547174
rect 294102 546618 294134 547174
rect 293514 511174 294134 546618
rect 293514 510618 293546 511174
rect 294102 510618 294134 511174
rect 293514 475174 294134 510618
rect 293514 474618 293546 475174
rect 294102 474618 294134 475174
rect 293514 439174 294134 474618
rect 293514 438618 293546 439174
rect 294102 438618 294134 439174
rect 293514 403174 294134 438618
rect 293514 402618 293546 403174
rect 294102 402618 294134 403174
rect 293514 367174 294134 402618
rect 293514 366618 293546 367174
rect 294102 366618 294134 367174
rect 293514 331174 294134 366618
rect 293514 330618 293546 331174
rect 294102 330618 294134 331174
rect 289794 326898 289826 327454
rect 290382 326898 290414 327454
rect 289794 291454 290414 326898
rect 292688 327454 293008 327486
rect 292688 327218 292730 327454
rect 292966 327218 293008 327454
rect 292688 327134 293008 327218
rect 292688 326898 292730 327134
rect 292966 326898 293008 327134
rect 292688 326866 293008 326898
rect 293514 295174 294134 330618
rect 293514 294618 293546 295174
rect 294102 294618 294134 295174
rect 289794 290898 289826 291454
rect 290382 290898 290414 291454
rect 289794 255454 290414 290898
rect 292688 291454 293008 291486
rect 292688 291218 292730 291454
rect 292966 291218 293008 291454
rect 292688 291134 293008 291218
rect 292688 290898 292730 291134
rect 292966 290898 293008 291134
rect 292688 290866 293008 290898
rect 293514 259174 294134 294618
rect 293514 258618 293546 259174
rect 294102 258618 294134 259174
rect 289794 254898 289826 255454
rect 290382 254898 290414 255454
rect 289794 219454 290414 254898
rect 292688 255454 293008 255486
rect 292688 255218 292730 255454
rect 292966 255218 293008 255454
rect 292688 255134 293008 255218
rect 292688 254898 292730 255134
rect 292966 254898 293008 255134
rect 292688 254866 293008 254898
rect 293514 223174 294134 258618
rect 293514 222618 293546 223174
rect 294102 222618 294134 223174
rect 289794 218898 289826 219454
rect 290382 218898 290414 219454
rect 289794 183454 290414 218898
rect 292688 219454 293008 219486
rect 292688 219218 292730 219454
rect 292966 219218 293008 219454
rect 292688 219134 293008 219218
rect 292688 218898 292730 219134
rect 292966 218898 293008 219134
rect 292688 218866 293008 218898
rect 293514 187174 294134 222618
rect 293514 186618 293546 187174
rect 294102 186618 294134 187174
rect 289794 182898 289826 183454
rect 290382 182898 290414 183454
rect 289794 147454 290414 182898
rect 292688 183454 293008 183486
rect 292688 183218 292730 183454
rect 292966 183218 293008 183454
rect 292688 183134 293008 183218
rect 292688 182898 292730 183134
rect 292966 182898 293008 183134
rect 292688 182866 293008 182898
rect 293514 151174 294134 186618
rect 293514 150618 293546 151174
rect 294102 150618 294134 151174
rect 289794 146898 289826 147454
rect 290382 146898 290414 147454
rect 289794 111454 290414 146898
rect 292688 147454 293008 147486
rect 292688 147218 292730 147454
rect 292966 147218 293008 147454
rect 292688 147134 293008 147218
rect 292688 146898 292730 147134
rect 292966 146898 293008 147134
rect 292688 146866 293008 146898
rect 293514 115174 294134 150618
rect 293514 114618 293546 115174
rect 294102 114618 294134 115174
rect 289794 110898 289826 111454
rect 290382 110898 290414 111454
rect 289794 75454 290414 110898
rect 292688 111454 293008 111486
rect 292688 111218 292730 111454
rect 292966 111218 293008 111454
rect 292688 111134 293008 111218
rect 292688 110898 292730 111134
rect 292966 110898 293008 111134
rect 292688 110866 293008 110898
rect 293514 79174 294134 114618
rect 293514 78618 293546 79174
rect 294102 78618 294134 79174
rect 289794 74898 289826 75454
rect 290382 74898 290414 75454
rect 289794 39454 290414 74898
rect 292688 75454 293008 75486
rect 292688 75218 292730 75454
rect 292966 75218 293008 75454
rect 292688 75134 293008 75218
rect 292688 74898 292730 75134
rect 292966 74898 293008 75134
rect 292688 74866 293008 74898
rect 293514 43174 294134 78618
rect 293514 42618 293546 43174
rect 294102 42618 294134 43174
rect 289794 38898 289826 39454
rect 290382 38898 290414 39454
rect 289794 3454 290414 38898
rect 292688 39454 293008 39486
rect 292688 39218 292730 39454
rect 292966 39218 293008 39454
rect 292688 39134 293008 39218
rect 292688 38898 292730 39134
rect 292966 38898 293008 39134
rect 292688 38866 293008 38898
rect 289794 2898 289826 3454
rect 290382 2898 290414 3454
rect 289794 -346 290414 2898
rect 289794 -902 289826 -346
rect 290382 -902 290414 -346
rect 289794 -7654 290414 -902
rect 293514 7174 294134 42618
rect 293514 6618 293546 7174
rect 294102 6618 294134 7174
rect 293514 -1306 294134 6618
rect 293514 -1862 293546 -1306
rect 294102 -1862 294134 -1306
rect 293514 -7654 294134 -1862
rect 297234 706758 297854 711590
rect 297234 706202 297266 706758
rect 297822 706202 297854 706758
rect 297234 694894 297854 706202
rect 297234 694338 297266 694894
rect 297822 694338 297854 694894
rect 297234 658894 297854 694338
rect 297234 658338 297266 658894
rect 297822 658338 297854 658894
rect 297234 622894 297854 658338
rect 297234 622338 297266 622894
rect 297822 622338 297854 622894
rect 297234 586894 297854 622338
rect 297234 586338 297266 586894
rect 297822 586338 297854 586894
rect 297234 550894 297854 586338
rect 297234 550338 297266 550894
rect 297822 550338 297854 550894
rect 297234 514894 297854 550338
rect 297234 514338 297266 514894
rect 297822 514338 297854 514894
rect 297234 478894 297854 514338
rect 297234 478338 297266 478894
rect 297822 478338 297854 478894
rect 297234 442894 297854 478338
rect 297234 442338 297266 442894
rect 297822 442338 297854 442894
rect 297234 406894 297854 442338
rect 297234 406338 297266 406894
rect 297822 406338 297854 406894
rect 297234 370894 297854 406338
rect 297234 370338 297266 370894
rect 297822 370338 297854 370894
rect 297234 334894 297854 370338
rect 297234 334338 297266 334894
rect 297822 334338 297854 334894
rect 297234 298894 297854 334338
rect 297234 298338 297266 298894
rect 297822 298338 297854 298894
rect 297234 262894 297854 298338
rect 297234 262338 297266 262894
rect 297822 262338 297854 262894
rect 297234 226894 297854 262338
rect 297234 226338 297266 226894
rect 297822 226338 297854 226894
rect 297234 190894 297854 226338
rect 297234 190338 297266 190894
rect 297822 190338 297854 190894
rect 297234 154894 297854 190338
rect 297234 154338 297266 154894
rect 297822 154338 297854 154894
rect 297234 118894 297854 154338
rect 297234 118338 297266 118894
rect 297822 118338 297854 118894
rect 297234 82894 297854 118338
rect 297234 82338 297266 82894
rect 297822 82338 297854 82894
rect 297234 46894 297854 82338
rect 297234 46338 297266 46894
rect 297822 46338 297854 46894
rect 297234 10894 297854 46338
rect 297234 10338 297266 10894
rect 297822 10338 297854 10894
rect 297234 -2266 297854 10338
rect 297234 -2822 297266 -2266
rect 297822 -2822 297854 -2266
rect 297234 -7654 297854 -2822
rect 300954 707718 301574 711590
rect 300954 707162 300986 707718
rect 301542 707162 301574 707718
rect 300954 698614 301574 707162
rect 300954 698058 300986 698614
rect 301542 698058 301574 698614
rect 300954 662614 301574 698058
rect 300954 662058 300986 662614
rect 301542 662058 301574 662614
rect 300954 626614 301574 662058
rect 300954 626058 300986 626614
rect 301542 626058 301574 626614
rect 300954 590614 301574 626058
rect 300954 590058 300986 590614
rect 301542 590058 301574 590614
rect 300954 554614 301574 590058
rect 300954 554058 300986 554614
rect 301542 554058 301574 554614
rect 300954 518614 301574 554058
rect 300954 518058 300986 518614
rect 301542 518058 301574 518614
rect 300954 482614 301574 518058
rect 300954 482058 300986 482614
rect 301542 482058 301574 482614
rect 300954 446614 301574 482058
rect 300954 446058 300986 446614
rect 301542 446058 301574 446614
rect 300954 410614 301574 446058
rect 300954 410058 300986 410614
rect 301542 410058 301574 410614
rect 300954 374614 301574 410058
rect 300954 374058 300986 374614
rect 301542 374058 301574 374614
rect 300954 338614 301574 374058
rect 300954 338058 300986 338614
rect 301542 338058 301574 338614
rect 300954 302614 301574 338058
rect 300954 302058 300986 302614
rect 301542 302058 301574 302614
rect 300954 266614 301574 302058
rect 300954 266058 300986 266614
rect 301542 266058 301574 266614
rect 300954 230614 301574 266058
rect 300954 230058 300986 230614
rect 301542 230058 301574 230614
rect 300954 194614 301574 230058
rect 300954 194058 300986 194614
rect 301542 194058 301574 194614
rect 300954 158614 301574 194058
rect 300954 158058 300986 158614
rect 301542 158058 301574 158614
rect 300954 122614 301574 158058
rect 300954 122058 300986 122614
rect 301542 122058 301574 122614
rect 300954 86614 301574 122058
rect 300954 86058 300986 86614
rect 301542 86058 301574 86614
rect 300954 50614 301574 86058
rect 300954 50058 300986 50614
rect 301542 50058 301574 50614
rect 300954 14614 301574 50058
rect 300954 14058 300986 14614
rect 301542 14058 301574 14614
rect 300954 -3226 301574 14058
rect 300954 -3782 300986 -3226
rect 301542 -3782 301574 -3226
rect 300954 -7654 301574 -3782
rect 304674 708678 305294 711590
rect 304674 708122 304706 708678
rect 305262 708122 305294 708678
rect 304674 666334 305294 708122
rect 304674 665778 304706 666334
rect 305262 665778 305294 666334
rect 304674 630334 305294 665778
rect 304674 629778 304706 630334
rect 305262 629778 305294 630334
rect 304674 594334 305294 629778
rect 304674 593778 304706 594334
rect 305262 593778 305294 594334
rect 304674 558334 305294 593778
rect 304674 557778 304706 558334
rect 305262 557778 305294 558334
rect 304674 522334 305294 557778
rect 304674 521778 304706 522334
rect 305262 521778 305294 522334
rect 304674 486334 305294 521778
rect 304674 485778 304706 486334
rect 305262 485778 305294 486334
rect 304674 450334 305294 485778
rect 304674 449778 304706 450334
rect 305262 449778 305294 450334
rect 304674 414334 305294 449778
rect 304674 413778 304706 414334
rect 305262 413778 305294 414334
rect 304674 378334 305294 413778
rect 304674 377778 304706 378334
rect 305262 377778 305294 378334
rect 304674 342334 305294 377778
rect 308394 709638 309014 711590
rect 308394 709082 308426 709638
rect 308982 709082 309014 709638
rect 308394 670054 309014 709082
rect 308394 669498 308426 670054
rect 308982 669498 309014 670054
rect 308394 634054 309014 669498
rect 308394 633498 308426 634054
rect 308982 633498 309014 634054
rect 308394 598054 309014 633498
rect 308394 597498 308426 598054
rect 308982 597498 309014 598054
rect 308394 562054 309014 597498
rect 308394 561498 308426 562054
rect 308982 561498 309014 562054
rect 308394 526054 309014 561498
rect 308394 525498 308426 526054
rect 308982 525498 309014 526054
rect 308394 490054 309014 525498
rect 308394 489498 308426 490054
rect 308982 489498 309014 490054
rect 308394 454054 309014 489498
rect 308394 453498 308426 454054
rect 308982 453498 309014 454054
rect 308394 418054 309014 453498
rect 308394 417498 308426 418054
rect 308982 417498 309014 418054
rect 308394 382054 309014 417498
rect 308394 381498 308426 382054
rect 308982 381498 309014 382054
rect 308394 354900 309014 381498
rect 312114 710598 312734 711590
rect 312114 710042 312146 710598
rect 312702 710042 312734 710598
rect 312114 673774 312734 710042
rect 312114 673218 312146 673774
rect 312702 673218 312734 673774
rect 312114 637774 312734 673218
rect 312114 637218 312146 637774
rect 312702 637218 312734 637774
rect 312114 601774 312734 637218
rect 312114 601218 312146 601774
rect 312702 601218 312734 601774
rect 312114 565774 312734 601218
rect 312114 565218 312146 565774
rect 312702 565218 312734 565774
rect 312114 529774 312734 565218
rect 312114 529218 312146 529774
rect 312702 529218 312734 529774
rect 312114 493774 312734 529218
rect 312114 493218 312146 493774
rect 312702 493218 312734 493774
rect 312114 457774 312734 493218
rect 312114 457218 312146 457774
rect 312702 457218 312734 457774
rect 312114 421774 312734 457218
rect 312114 421218 312146 421774
rect 312702 421218 312734 421774
rect 312114 385774 312734 421218
rect 312114 385218 312146 385774
rect 312702 385218 312734 385774
rect 304674 341778 304706 342334
rect 305262 341778 305294 342334
rect 304674 306334 305294 341778
rect 312114 349774 312734 385218
rect 312114 349218 312146 349774
rect 312702 349218 312734 349774
rect 308048 331174 308368 331206
rect 308048 330938 308090 331174
rect 308326 330938 308368 331174
rect 308048 330854 308368 330938
rect 308048 330618 308090 330854
rect 308326 330618 308368 330854
rect 308048 330586 308368 330618
rect 304674 305778 304706 306334
rect 305262 305778 305294 306334
rect 304674 270334 305294 305778
rect 312114 313774 312734 349218
rect 312114 313218 312146 313774
rect 312702 313218 312734 313774
rect 308048 295174 308368 295206
rect 308048 294938 308090 295174
rect 308326 294938 308368 295174
rect 308048 294854 308368 294938
rect 308048 294618 308090 294854
rect 308326 294618 308368 294854
rect 308048 294586 308368 294618
rect 304674 269778 304706 270334
rect 305262 269778 305294 270334
rect 304674 234334 305294 269778
rect 312114 277774 312734 313218
rect 312114 277218 312146 277774
rect 312702 277218 312734 277774
rect 308048 259174 308368 259206
rect 308048 258938 308090 259174
rect 308326 258938 308368 259174
rect 308048 258854 308368 258938
rect 308048 258618 308090 258854
rect 308326 258618 308368 258854
rect 308048 258586 308368 258618
rect 304674 233778 304706 234334
rect 305262 233778 305294 234334
rect 304674 198334 305294 233778
rect 312114 241774 312734 277218
rect 312114 241218 312146 241774
rect 312702 241218 312734 241774
rect 308048 223174 308368 223206
rect 308048 222938 308090 223174
rect 308326 222938 308368 223174
rect 308048 222854 308368 222938
rect 308048 222618 308090 222854
rect 308326 222618 308368 222854
rect 308048 222586 308368 222618
rect 304674 197778 304706 198334
rect 305262 197778 305294 198334
rect 304674 162334 305294 197778
rect 312114 205774 312734 241218
rect 312114 205218 312146 205774
rect 312702 205218 312734 205774
rect 308048 187174 308368 187206
rect 308048 186938 308090 187174
rect 308326 186938 308368 187174
rect 308048 186854 308368 186938
rect 308048 186618 308090 186854
rect 308326 186618 308368 186854
rect 308048 186586 308368 186618
rect 304674 161778 304706 162334
rect 305262 161778 305294 162334
rect 304674 126334 305294 161778
rect 312114 169774 312734 205218
rect 312114 169218 312146 169774
rect 312702 169218 312734 169774
rect 308048 151174 308368 151206
rect 308048 150938 308090 151174
rect 308326 150938 308368 151174
rect 308048 150854 308368 150938
rect 308048 150618 308090 150854
rect 308326 150618 308368 150854
rect 308048 150586 308368 150618
rect 304674 125778 304706 126334
rect 305262 125778 305294 126334
rect 304674 90334 305294 125778
rect 312114 133774 312734 169218
rect 312114 133218 312146 133774
rect 312702 133218 312734 133774
rect 308048 115174 308368 115206
rect 308048 114938 308090 115174
rect 308326 114938 308368 115174
rect 308048 114854 308368 114938
rect 308048 114618 308090 114854
rect 308326 114618 308368 114854
rect 308048 114586 308368 114618
rect 304674 89778 304706 90334
rect 305262 89778 305294 90334
rect 304674 54334 305294 89778
rect 312114 97774 312734 133218
rect 312114 97218 312146 97774
rect 312702 97218 312734 97774
rect 308048 79174 308368 79206
rect 308048 78938 308090 79174
rect 308326 78938 308368 79174
rect 308048 78854 308368 78938
rect 308048 78618 308090 78854
rect 308326 78618 308368 78854
rect 308048 78586 308368 78618
rect 304674 53778 304706 54334
rect 305262 53778 305294 54334
rect 304674 18334 305294 53778
rect 312114 61774 312734 97218
rect 312114 61218 312146 61774
rect 312702 61218 312734 61774
rect 308048 43174 308368 43206
rect 308048 42938 308090 43174
rect 308326 42938 308368 43174
rect 308048 42854 308368 42938
rect 308048 42618 308090 42854
rect 308326 42618 308368 42854
rect 308048 42586 308368 42618
rect 304674 17778 304706 18334
rect 305262 17778 305294 18334
rect 304674 -4186 305294 17778
rect 312114 25774 312734 61218
rect 312114 25218 312146 25774
rect 312702 25218 312734 25774
rect 308048 7174 308368 7206
rect 308048 6938 308090 7174
rect 308326 6938 308368 7174
rect 308048 6854 308368 6938
rect 308048 6618 308090 6854
rect 308326 6618 308368 6854
rect 308048 6586 308368 6618
rect 304674 -4742 304706 -4186
rect 305262 -4742 305294 -4186
rect 304674 -7654 305294 -4742
rect 312114 -6106 312734 25218
rect 312114 -6662 312146 -6106
rect 312702 -6662 312734 -6106
rect 312114 -7654 312734 -6662
rect 315834 711558 316454 711590
rect 315834 711002 315866 711558
rect 316422 711002 316454 711558
rect 315834 677494 316454 711002
rect 315834 676938 315866 677494
rect 316422 676938 316454 677494
rect 315834 641494 316454 676938
rect 315834 640938 315866 641494
rect 316422 640938 316454 641494
rect 315834 605494 316454 640938
rect 315834 604938 315866 605494
rect 316422 604938 316454 605494
rect 315834 569494 316454 604938
rect 315834 568938 315866 569494
rect 316422 568938 316454 569494
rect 315834 533494 316454 568938
rect 315834 532938 315866 533494
rect 316422 532938 316454 533494
rect 315834 497494 316454 532938
rect 315834 496938 315866 497494
rect 316422 496938 316454 497494
rect 315834 461494 316454 496938
rect 315834 460938 315866 461494
rect 316422 460938 316454 461494
rect 315834 425494 316454 460938
rect 315834 424938 315866 425494
rect 316422 424938 316454 425494
rect 315834 389494 316454 424938
rect 315834 388938 315866 389494
rect 316422 388938 316454 389494
rect 315834 353494 316454 388938
rect 315834 352938 315866 353494
rect 316422 352938 316454 353494
rect 315834 317494 316454 352938
rect 325794 704838 326414 711590
rect 325794 704282 325826 704838
rect 326382 704282 326414 704838
rect 325794 687454 326414 704282
rect 325794 686898 325826 687454
rect 326382 686898 326414 687454
rect 325794 651454 326414 686898
rect 325794 650898 325826 651454
rect 326382 650898 326414 651454
rect 325794 615454 326414 650898
rect 325794 614898 325826 615454
rect 326382 614898 326414 615454
rect 325794 579454 326414 614898
rect 325794 578898 325826 579454
rect 326382 578898 326414 579454
rect 325794 543454 326414 578898
rect 325794 542898 325826 543454
rect 326382 542898 326414 543454
rect 325794 507454 326414 542898
rect 325794 506898 325826 507454
rect 326382 506898 326414 507454
rect 325794 471454 326414 506898
rect 325794 470898 325826 471454
rect 326382 470898 326414 471454
rect 325794 435454 326414 470898
rect 325794 434898 325826 435454
rect 326382 434898 326414 435454
rect 325794 399454 326414 434898
rect 325794 398898 325826 399454
rect 326382 398898 326414 399454
rect 325794 363454 326414 398898
rect 325794 362898 325826 363454
rect 326382 362898 326414 363454
rect 323408 327454 323728 327486
rect 323408 327218 323450 327454
rect 323686 327218 323728 327454
rect 323408 327134 323728 327218
rect 323408 326898 323450 327134
rect 323686 326898 323728 327134
rect 323408 326866 323728 326898
rect 325794 327454 326414 362898
rect 325794 326898 325826 327454
rect 326382 326898 326414 327454
rect 315834 316938 315866 317494
rect 316422 316938 316454 317494
rect 315834 281494 316454 316938
rect 323408 291454 323728 291486
rect 323408 291218 323450 291454
rect 323686 291218 323728 291454
rect 323408 291134 323728 291218
rect 323408 290898 323450 291134
rect 323686 290898 323728 291134
rect 323408 290866 323728 290898
rect 325794 291454 326414 326898
rect 325794 290898 325826 291454
rect 326382 290898 326414 291454
rect 315834 280938 315866 281494
rect 316422 280938 316454 281494
rect 315834 245494 316454 280938
rect 323408 255454 323728 255486
rect 323408 255218 323450 255454
rect 323686 255218 323728 255454
rect 323408 255134 323728 255218
rect 323408 254898 323450 255134
rect 323686 254898 323728 255134
rect 323408 254866 323728 254898
rect 325794 255454 326414 290898
rect 325794 254898 325826 255454
rect 326382 254898 326414 255454
rect 315834 244938 315866 245494
rect 316422 244938 316454 245494
rect 315834 209494 316454 244938
rect 323408 219454 323728 219486
rect 323408 219218 323450 219454
rect 323686 219218 323728 219454
rect 323408 219134 323728 219218
rect 323408 218898 323450 219134
rect 323686 218898 323728 219134
rect 323408 218866 323728 218898
rect 325794 219454 326414 254898
rect 325794 218898 325826 219454
rect 326382 218898 326414 219454
rect 315834 208938 315866 209494
rect 316422 208938 316454 209494
rect 315834 173494 316454 208938
rect 323408 183454 323728 183486
rect 323408 183218 323450 183454
rect 323686 183218 323728 183454
rect 323408 183134 323728 183218
rect 323408 182898 323450 183134
rect 323686 182898 323728 183134
rect 323408 182866 323728 182898
rect 325794 183454 326414 218898
rect 325794 182898 325826 183454
rect 326382 182898 326414 183454
rect 315834 172938 315866 173494
rect 316422 172938 316454 173494
rect 315834 137494 316454 172938
rect 323408 147454 323728 147486
rect 323408 147218 323450 147454
rect 323686 147218 323728 147454
rect 323408 147134 323728 147218
rect 323408 146898 323450 147134
rect 323686 146898 323728 147134
rect 323408 146866 323728 146898
rect 325794 147454 326414 182898
rect 325794 146898 325826 147454
rect 326382 146898 326414 147454
rect 315834 136938 315866 137494
rect 316422 136938 316454 137494
rect 315834 101494 316454 136938
rect 323408 111454 323728 111486
rect 323408 111218 323450 111454
rect 323686 111218 323728 111454
rect 323408 111134 323728 111218
rect 323408 110898 323450 111134
rect 323686 110898 323728 111134
rect 323408 110866 323728 110898
rect 325794 111454 326414 146898
rect 325794 110898 325826 111454
rect 326382 110898 326414 111454
rect 315834 100938 315866 101494
rect 316422 100938 316454 101494
rect 315834 65494 316454 100938
rect 323408 75454 323728 75486
rect 323408 75218 323450 75454
rect 323686 75218 323728 75454
rect 323408 75134 323728 75218
rect 323408 74898 323450 75134
rect 323686 74898 323728 75134
rect 323408 74866 323728 74898
rect 325794 75454 326414 110898
rect 325794 74898 325826 75454
rect 326382 74898 326414 75454
rect 315834 64938 315866 65494
rect 316422 64938 316454 65494
rect 315834 29494 316454 64938
rect 323408 39454 323728 39486
rect 323408 39218 323450 39454
rect 323686 39218 323728 39454
rect 323408 39134 323728 39218
rect 323408 38898 323450 39134
rect 323686 38898 323728 39134
rect 323408 38866 323728 38898
rect 325794 39454 326414 74898
rect 325794 38898 325826 39454
rect 326382 38898 326414 39454
rect 315834 28938 315866 29494
rect 316422 28938 316454 29494
rect 315834 -7066 316454 28938
rect 315834 -7622 315866 -7066
rect 316422 -7622 316454 -7066
rect 315834 -7654 316454 -7622
rect 325794 3454 326414 38898
rect 325794 2898 325826 3454
rect 326382 2898 326414 3454
rect 325794 -346 326414 2898
rect 325794 -902 325826 -346
rect 326382 -902 326414 -346
rect 325794 -7654 326414 -902
rect 329514 705798 330134 711590
rect 329514 705242 329546 705798
rect 330102 705242 330134 705798
rect 329514 691174 330134 705242
rect 329514 690618 329546 691174
rect 330102 690618 330134 691174
rect 329514 655174 330134 690618
rect 329514 654618 329546 655174
rect 330102 654618 330134 655174
rect 329514 619174 330134 654618
rect 329514 618618 329546 619174
rect 330102 618618 330134 619174
rect 329514 583174 330134 618618
rect 329514 582618 329546 583174
rect 330102 582618 330134 583174
rect 329514 547174 330134 582618
rect 329514 546618 329546 547174
rect 330102 546618 330134 547174
rect 329514 511174 330134 546618
rect 329514 510618 329546 511174
rect 330102 510618 330134 511174
rect 329514 475174 330134 510618
rect 329514 474618 329546 475174
rect 330102 474618 330134 475174
rect 329514 439174 330134 474618
rect 329514 438618 329546 439174
rect 330102 438618 330134 439174
rect 329514 403174 330134 438618
rect 329514 402618 329546 403174
rect 330102 402618 330134 403174
rect 329514 367174 330134 402618
rect 329514 366618 329546 367174
rect 330102 366618 330134 367174
rect 329514 331174 330134 366618
rect 329514 330618 329546 331174
rect 330102 330618 330134 331174
rect 329514 295174 330134 330618
rect 329514 294618 329546 295174
rect 330102 294618 330134 295174
rect 329514 259174 330134 294618
rect 329514 258618 329546 259174
rect 330102 258618 330134 259174
rect 329514 223174 330134 258618
rect 329514 222618 329546 223174
rect 330102 222618 330134 223174
rect 329514 187174 330134 222618
rect 329514 186618 329546 187174
rect 330102 186618 330134 187174
rect 329514 151174 330134 186618
rect 329514 150618 329546 151174
rect 330102 150618 330134 151174
rect 329514 115174 330134 150618
rect 329514 114618 329546 115174
rect 330102 114618 330134 115174
rect 329514 79174 330134 114618
rect 329514 78618 329546 79174
rect 330102 78618 330134 79174
rect 329514 43174 330134 78618
rect 329514 42618 329546 43174
rect 330102 42618 330134 43174
rect 329514 7174 330134 42618
rect 329514 6618 329546 7174
rect 330102 6618 330134 7174
rect 329514 -1306 330134 6618
rect 329514 -1862 329546 -1306
rect 330102 -1862 330134 -1306
rect 329514 -7654 330134 -1862
rect 333234 706758 333854 711590
rect 333234 706202 333266 706758
rect 333822 706202 333854 706758
rect 333234 694894 333854 706202
rect 333234 694338 333266 694894
rect 333822 694338 333854 694894
rect 333234 658894 333854 694338
rect 333234 658338 333266 658894
rect 333822 658338 333854 658894
rect 333234 622894 333854 658338
rect 333234 622338 333266 622894
rect 333822 622338 333854 622894
rect 333234 586894 333854 622338
rect 333234 586338 333266 586894
rect 333822 586338 333854 586894
rect 333234 550894 333854 586338
rect 333234 550338 333266 550894
rect 333822 550338 333854 550894
rect 333234 514894 333854 550338
rect 333234 514338 333266 514894
rect 333822 514338 333854 514894
rect 333234 478894 333854 514338
rect 333234 478338 333266 478894
rect 333822 478338 333854 478894
rect 333234 442894 333854 478338
rect 333234 442338 333266 442894
rect 333822 442338 333854 442894
rect 333234 406894 333854 442338
rect 333234 406338 333266 406894
rect 333822 406338 333854 406894
rect 333234 370894 333854 406338
rect 333234 370338 333266 370894
rect 333822 370338 333854 370894
rect 333234 334894 333854 370338
rect 333234 334338 333266 334894
rect 333822 334338 333854 334894
rect 333234 298894 333854 334338
rect 333234 298338 333266 298894
rect 333822 298338 333854 298894
rect 333234 262894 333854 298338
rect 333234 262338 333266 262894
rect 333822 262338 333854 262894
rect 333234 226894 333854 262338
rect 333234 226338 333266 226894
rect 333822 226338 333854 226894
rect 333234 190894 333854 226338
rect 333234 190338 333266 190894
rect 333822 190338 333854 190894
rect 333234 154894 333854 190338
rect 333234 154338 333266 154894
rect 333822 154338 333854 154894
rect 333234 118894 333854 154338
rect 333234 118338 333266 118894
rect 333822 118338 333854 118894
rect 333234 82894 333854 118338
rect 333234 82338 333266 82894
rect 333822 82338 333854 82894
rect 333234 46894 333854 82338
rect 333234 46338 333266 46894
rect 333822 46338 333854 46894
rect 333234 10894 333854 46338
rect 333234 10338 333266 10894
rect 333822 10338 333854 10894
rect 333234 -2266 333854 10338
rect 333234 -2822 333266 -2266
rect 333822 -2822 333854 -2266
rect 333234 -7654 333854 -2822
rect 336954 707718 337574 711590
rect 336954 707162 336986 707718
rect 337542 707162 337574 707718
rect 336954 698614 337574 707162
rect 336954 698058 336986 698614
rect 337542 698058 337574 698614
rect 336954 662614 337574 698058
rect 336954 662058 336986 662614
rect 337542 662058 337574 662614
rect 336954 626614 337574 662058
rect 336954 626058 336986 626614
rect 337542 626058 337574 626614
rect 336954 590614 337574 626058
rect 336954 590058 336986 590614
rect 337542 590058 337574 590614
rect 336954 554614 337574 590058
rect 336954 554058 336986 554614
rect 337542 554058 337574 554614
rect 336954 518614 337574 554058
rect 336954 518058 336986 518614
rect 337542 518058 337574 518614
rect 336954 482614 337574 518058
rect 336954 482058 336986 482614
rect 337542 482058 337574 482614
rect 336954 446614 337574 482058
rect 336954 446058 336986 446614
rect 337542 446058 337574 446614
rect 336954 410614 337574 446058
rect 336954 410058 336986 410614
rect 337542 410058 337574 410614
rect 336954 374614 337574 410058
rect 336954 374058 336986 374614
rect 337542 374058 337574 374614
rect 336954 338614 337574 374058
rect 336954 338058 336986 338614
rect 337542 338058 337574 338614
rect 336954 302614 337574 338058
rect 340674 708678 341294 711590
rect 340674 708122 340706 708678
rect 341262 708122 341294 708678
rect 340674 666334 341294 708122
rect 340674 665778 340706 666334
rect 341262 665778 341294 666334
rect 340674 630334 341294 665778
rect 340674 629778 340706 630334
rect 341262 629778 341294 630334
rect 340674 594334 341294 629778
rect 340674 593778 340706 594334
rect 341262 593778 341294 594334
rect 340674 558334 341294 593778
rect 340674 557778 340706 558334
rect 341262 557778 341294 558334
rect 340674 522334 341294 557778
rect 340674 521778 340706 522334
rect 341262 521778 341294 522334
rect 340674 486334 341294 521778
rect 340674 485778 340706 486334
rect 341262 485778 341294 486334
rect 340674 450334 341294 485778
rect 340674 449778 340706 450334
rect 341262 449778 341294 450334
rect 340674 414334 341294 449778
rect 340674 413778 340706 414334
rect 341262 413778 341294 414334
rect 340674 378334 341294 413778
rect 340674 377778 340706 378334
rect 341262 377778 341294 378334
rect 340674 342334 341294 377778
rect 340674 341778 340706 342334
rect 341262 341778 341294 342334
rect 338768 331174 339088 331206
rect 338768 330938 338810 331174
rect 339046 330938 339088 331174
rect 338768 330854 339088 330938
rect 338768 330618 338810 330854
rect 339046 330618 339088 330854
rect 338768 330586 339088 330618
rect 336954 302058 336986 302614
rect 337542 302058 337574 302614
rect 336954 266614 337574 302058
rect 340674 306334 341294 341778
rect 340674 305778 340706 306334
rect 341262 305778 341294 306334
rect 338768 295174 339088 295206
rect 338768 294938 338810 295174
rect 339046 294938 339088 295174
rect 338768 294854 339088 294938
rect 338768 294618 338810 294854
rect 339046 294618 339088 294854
rect 338768 294586 339088 294618
rect 336954 266058 336986 266614
rect 337542 266058 337574 266614
rect 336954 230614 337574 266058
rect 340674 270334 341294 305778
rect 340674 269778 340706 270334
rect 341262 269778 341294 270334
rect 338768 259174 339088 259206
rect 338768 258938 338810 259174
rect 339046 258938 339088 259174
rect 338768 258854 339088 258938
rect 338768 258618 338810 258854
rect 339046 258618 339088 258854
rect 338768 258586 339088 258618
rect 336954 230058 336986 230614
rect 337542 230058 337574 230614
rect 336954 194614 337574 230058
rect 340674 234334 341294 269778
rect 340674 233778 340706 234334
rect 341262 233778 341294 234334
rect 338768 223174 339088 223206
rect 338768 222938 338810 223174
rect 339046 222938 339088 223174
rect 338768 222854 339088 222938
rect 338768 222618 338810 222854
rect 339046 222618 339088 222854
rect 338768 222586 339088 222618
rect 336954 194058 336986 194614
rect 337542 194058 337574 194614
rect 336954 158614 337574 194058
rect 340674 198334 341294 233778
rect 340674 197778 340706 198334
rect 341262 197778 341294 198334
rect 338768 187174 339088 187206
rect 338768 186938 338810 187174
rect 339046 186938 339088 187174
rect 338768 186854 339088 186938
rect 338768 186618 338810 186854
rect 339046 186618 339088 186854
rect 338768 186586 339088 186618
rect 336954 158058 336986 158614
rect 337542 158058 337574 158614
rect 336954 122614 337574 158058
rect 340674 162334 341294 197778
rect 340674 161778 340706 162334
rect 341262 161778 341294 162334
rect 338768 151174 339088 151206
rect 338768 150938 338810 151174
rect 339046 150938 339088 151174
rect 338768 150854 339088 150938
rect 338768 150618 338810 150854
rect 339046 150618 339088 150854
rect 338768 150586 339088 150618
rect 336954 122058 336986 122614
rect 337542 122058 337574 122614
rect 336954 86614 337574 122058
rect 340674 126334 341294 161778
rect 340674 125778 340706 126334
rect 341262 125778 341294 126334
rect 338768 115174 339088 115206
rect 338768 114938 338810 115174
rect 339046 114938 339088 115174
rect 338768 114854 339088 114938
rect 338768 114618 338810 114854
rect 339046 114618 339088 114854
rect 338768 114586 339088 114618
rect 336954 86058 336986 86614
rect 337542 86058 337574 86614
rect 336954 50614 337574 86058
rect 340674 90334 341294 125778
rect 340674 89778 340706 90334
rect 341262 89778 341294 90334
rect 338768 79174 339088 79206
rect 338768 78938 338810 79174
rect 339046 78938 339088 79174
rect 338768 78854 339088 78938
rect 338768 78618 338810 78854
rect 339046 78618 339088 78854
rect 338768 78586 339088 78618
rect 336954 50058 336986 50614
rect 337542 50058 337574 50614
rect 336954 14614 337574 50058
rect 340674 54334 341294 89778
rect 340674 53778 340706 54334
rect 341262 53778 341294 54334
rect 338768 43174 339088 43206
rect 338768 42938 338810 43174
rect 339046 42938 339088 43174
rect 338768 42854 339088 42938
rect 338768 42618 338810 42854
rect 339046 42618 339088 42854
rect 338768 42586 339088 42618
rect 336954 14058 336986 14614
rect 337542 14058 337574 14614
rect 336954 -3226 337574 14058
rect 340674 18334 341294 53778
rect 340674 17778 340706 18334
rect 341262 17778 341294 18334
rect 338768 7174 339088 7206
rect 338768 6938 338810 7174
rect 339046 6938 339088 7174
rect 338768 6854 339088 6938
rect 338768 6618 338810 6854
rect 339046 6618 339088 6854
rect 338768 6586 339088 6618
rect 336954 -3782 336986 -3226
rect 337542 -3782 337574 -3226
rect 336954 -7654 337574 -3782
rect 340674 -4186 341294 17778
rect 340674 -4742 340706 -4186
rect 341262 -4742 341294 -4186
rect 340674 -7654 341294 -4742
rect 344394 709638 345014 711590
rect 344394 709082 344426 709638
rect 344982 709082 345014 709638
rect 344394 670054 345014 709082
rect 344394 669498 344426 670054
rect 344982 669498 345014 670054
rect 344394 634054 345014 669498
rect 344394 633498 344426 634054
rect 344982 633498 345014 634054
rect 344394 598054 345014 633498
rect 344394 597498 344426 598054
rect 344982 597498 345014 598054
rect 344394 562054 345014 597498
rect 344394 561498 344426 562054
rect 344982 561498 345014 562054
rect 344394 526054 345014 561498
rect 344394 525498 344426 526054
rect 344982 525498 345014 526054
rect 344394 490054 345014 525498
rect 344394 489498 344426 490054
rect 344982 489498 345014 490054
rect 344394 454054 345014 489498
rect 344394 453498 344426 454054
rect 344982 453498 345014 454054
rect 344394 418054 345014 453498
rect 344394 417498 344426 418054
rect 344982 417498 345014 418054
rect 344394 382054 345014 417498
rect 344394 381498 344426 382054
rect 344982 381498 345014 382054
rect 344394 346054 345014 381498
rect 344394 345498 344426 346054
rect 344982 345498 345014 346054
rect 344394 310054 345014 345498
rect 344394 309498 344426 310054
rect 344982 309498 345014 310054
rect 344394 274054 345014 309498
rect 344394 273498 344426 274054
rect 344982 273498 345014 274054
rect 344394 238054 345014 273498
rect 344394 237498 344426 238054
rect 344982 237498 345014 238054
rect 344394 202054 345014 237498
rect 344394 201498 344426 202054
rect 344982 201498 345014 202054
rect 344394 166054 345014 201498
rect 344394 165498 344426 166054
rect 344982 165498 345014 166054
rect 344394 130054 345014 165498
rect 344394 129498 344426 130054
rect 344982 129498 345014 130054
rect 344394 94054 345014 129498
rect 344394 93498 344426 94054
rect 344982 93498 345014 94054
rect 344394 58054 345014 93498
rect 344394 57498 344426 58054
rect 344982 57498 345014 58054
rect 344394 22054 345014 57498
rect 344394 21498 344426 22054
rect 344982 21498 345014 22054
rect 344394 -5146 345014 21498
rect 344394 -5702 344426 -5146
rect 344982 -5702 345014 -5146
rect 344394 -7654 345014 -5702
rect 348114 710598 348734 711590
rect 348114 710042 348146 710598
rect 348702 710042 348734 710598
rect 348114 673774 348734 710042
rect 348114 673218 348146 673774
rect 348702 673218 348734 673774
rect 348114 637774 348734 673218
rect 348114 637218 348146 637774
rect 348702 637218 348734 637774
rect 348114 601774 348734 637218
rect 348114 601218 348146 601774
rect 348702 601218 348734 601774
rect 348114 565774 348734 601218
rect 348114 565218 348146 565774
rect 348702 565218 348734 565774
rect 348114 529774 348734 565218
rect 348114 529218 348146 529774
rect 348702 529218 348734 529774
rect 348114 493774 348734 529218
rect 348114 493218 348146 493774
rect 348702 493218 348734 493774
rect 348114 457774 348734 493218
rect 348114 457218 348146 457774
rect 348702 457218 348734 457774
rect 348114 421774 348734 457218
rect 348114 421218 348146 421774
rect 348702 421218 348734 421774
rect 348114 385774 348734 421218
rect 348114 385218 348146 385774
rect 348702 385218 348734 385774
rect 348114 349774 348734 385218
rect 348114 349218 348146 349774
rect 348702 349218 348734 349774
rect 348114 313774 348734 349218
rect 348114 313218 348146 313774
rect 348702 313218 348734 313774
rect 348114 277774 348734 313218
rect 348114 277218 348146 277774
rect 348702 277218 348734 277774
rect 348114 241774 348734 277218
rect 348114 241218 348146 241774
rect 348702 241218 348734 241774
rect 348114 205774 348734 241218
rect 348114 205218 348146 205774
rect 348702 205218 348734 205774
rect 348114 169774 348734 205218
rect 348114 169218 348146 169774
rect 348702 169218 348734 169774
rect 348114 133774 348734 169218
rect 348114 133218 348146 133774
rect 348702 133218 348734 133774
rect 348114 97774 348734 133218
rect 348114 97218 348146 97774
rect 348702 97218 348734 97774
rect 348114 61774 348734 97218
rect 348114 61218 348146 61774
rect 348702 61218 348734 61774
rect 348114 25774 348734 61218
rect 348114 25218 348146 25774
rect 348702 25218 348734 25774
rect 348114 -6106 348734 25218
rect 348114 -6662 348146 -6106
rect 348702 -6662 348734 -6106
rect 348114 -7654 348734 -6662
rect 351834 711558 352454 711590
rect 351834 711002 351866 711558
rect 352422 711002 352454 711558
rect 351834 677494 352454 711002
rect 351834 676938 351866 677494
rect 352422 676938 352454 677494
rect 351834 641494 352454 676938
rect 351834 640938 351866 641494
rect 352422 640938 352454 641494
rect 351834 605494 352454 640938
rect 351834 604938 351866 605494
rect 352422 604938 352454 605494
rect 351834 569494 352454 604938
rect 351834 568938 351866 569494
rect 352422 568938 352454 569494
rect 351834 533494 352454 568938
rect 351834 532938 351866 533494
rect 352422 532938 352454 533494
rect 351834 497494 352454 532938
rect 351834 496938 351866 497494
rect 352422 496938 352454 497494
rect 351834 461494 352454 496938
rect 351834 460938 351866 461494
rect 352422 460938 352454 461494
rect 351834 425494 352454 460938
rect 351834 424938 351866 425494
rect 352422 424938 352454 425494
rect 351834 389494 352454 424938
rect 351834 388938 351866 389494
rect 352422 388938 352454 389494
rect 351834 353494 352454 388938
rect 351834 352938 351866 353494
rect 352422 352938 352454 353494
rect 351834 317494 352454 352938
rect 361794 704838 362414 711590
rect 361794 704282 361826 704838
rect 362382 704282 362414 704838
rect 361794 687454 362414 704282
rect 361794 686898 361826 687454
rect 362382 686898 362414 687454
rect 361794 651454 362414 686898
rect 361794 650898 361826 651454
rect 362382 650898 362414 651454
rect 361794 615454 362414 650898
rect 361794 614898 361826 615454
rect 362382 614898 362414 615454
rect 361794 579454 362414 614898
rect 361794 578898 361826 579454
rect 362382 578898 362414 579454
rect 361794 543454 362414 578898
rect 361794 542898 361826 543454
rect 362382 542898 362414 543454
rect 361794 507454 362414 542898
rect 361794 506898 361826 507454
rect 362382 506898 362414 507454
rect 361794 471454 362414 506898
rect 361794 470898 361826 471454
rect 362382 470898 362414 471454
rect 361794 435454 362414 470898
rect 361794 434898 361826 435454
rect 362382 434898 362414 435454
rect 361794 399454 362414 434898
rect 361794 398898 361826 399454
rect 362382 398898 362414 399454
rect 361794 363454 362414 398898
rect 361794 362898 361826 363454
rect 362382 362898 362414 363454
rect 354128 327454 354448 327486
rect 354128 327218 354170 327454
rect 354406 327218 354448 327454
rect 354128 327134 354448 327218
rect 354128 326898 354170 327134
rect 354406 326898 354448 327134
rect 354128 326866 354448 326898
rect 361794 327454 362414 362898
rect 361794 326898 361826 327454
rect 362382 326898 362414 327454
rect 351834 316938 351866 317494
rect 352422 316938 352454 317494
rect 351834 281494 352454 316938
rect 354128 291454 354448 291486
rect 354128 291218 354170 291454
rect 354406 291218 354448 291454
rect 354128 291134 354448 291218
rect 354128 290898 354170 291134
rect 354406 290898 354448 291134
rect 354128 290866 354448 290898
rect 361794 291454 362414 326898
rect 361794 290898 361826 291454
rect 362382 290898 362414 291454
rect 351834 280938 351866 281494
rect 352422 280938 352454 281494
rect 351834 245494 352454 280938
rect 354128 255454 354448 255486
rect 354128 255218 354170 255454
rect 354406 255218 354448 255454
rect 354128 255134 354448 255218
rect 354128 254898 354170 255134
rect 354406 254898 354448 255134
rect 354128 254866 354448 254898
rect 361794 255454 362414 290898
rect 361794 254898 361826 255454
rect 362382 254898 362414 255454
rect 351834 244938 351866 245494
rect 352422 244938 352454 245494
rect 351834 209494 352454 244938
rect 354128 219454 354448 219486
rect 354128 219218 354170 219454
rect 354406 219218 354448 219454
rect 354128 219134 354448 219218
rect 354128 218898 354170 219134
rect 354406 218898 354448 219134
rect 354128 218866 354448 218898
rect 361794 219454 362414 254898
rect 361794 218898 361826 219454
rect 362382 218898 362414 219454
rect 351834 208938 351866 209494
rect 352422 208938 352454 209494
rect 351834 173494 352454 208938
rect 354128 183454 354448 183486
rect 354128 183218 354170 183454
rect 354406 183218 354448 183454
rect 354128 183134 354448 183218
rect 354128 182898 354170 183134
rect 354406 182898 354448 183134
rect 354128 182866 354448 182898
rect 361794 183454 362414 218898
rect 361794 182898 361826 183454
rect 362382 182898 362414 183454
rect 351834 172938 351866 173494
rect 352422 172938 352454 173494
rect 351834 137494 352454 172938
rect 354128 147454 354448 147486
rect 354128 147218 354170 147454
rect 354406 147218 354448 147454
rect 354128 147134 354448 147218
rect 354128 146898 354170 147134
rect 354406 146898 354448 147134
rect 354128 146866 354448 146898
rect 361794 147454 362414 182898
rect 361794 146898 361826 147454
rect 362382 146898 362414 147454
rect 351834 136938 351866 137494
rect 352422 136938 352454 137494
rect 351834 101494 352454 136938
rect 354128 111454 354448 111486
rect 354128 111218 354170 111454
rect 354406 111218 354448 111454
rect 354128 111134 354448 111218
rect 354128 110898 354170 111134
rect 354406 110898 354448 111134
rect 354128 110866 354448 110898
rect 361794 111454 362414 146898
rect 361794 110898 361826 111454
rect 362382 110898 362414 111454
rect 351834 100938 351866 101494
rect 352422 100938 352454 101494
rect 351834 65494 352454 100938
rect 354128 75454 354448 75486
rect 354128 75218 354170 75454
rect 354406 75218 354448 75454
rect 354128 75134 354448 75218
rect 354128 74898 354170 75134
rect 354406 74898 354448 75134
rect 354128 74866 354448 74898
rect 361794 75454 362414 110898
rect 361794 74898 361826 75454
rect 362382 74898 362414 75454
rect 351834 64938 351866 65494
rect 352422 64938 352454 65494
rect 351834 29494 352454 64938
rect 354128 39454 354448 39486
rect 354128 39218 354170 39454
rect 354406 39218 354448 39454
rect 354128 39134 354448 39218
rect 354128 38898 354170 39134
rect 354406 38898 354448 39134
rect 354128 38866 354448 38898
rect 361794 39454 362414 74898
rect 361794 38898 361826 39454
rect 362382 38898 362414 39454
rect 351834 28938 351866 29494
rect 352422 28938 352454 29494
rect 351834 -7066 352454 28938
rect 351834 -7622 351866 -7066
rect 352422 -7622 352454 -7066
rect 351834 -7654 352454 -7622
rect 361794 3454 362414 38898
rect 361794 2898 361826 3454
rect 362382 2898 362414 3454
rect 361794 -346 362414 2898
rect 361794 -902 361826 -346
rect 362382 -902 362414 -346
rect 361794 -7654 362414 -902
rect 365514 705798 366134 711590
rect 365514 705242 365546 705798
rect 366102 705242 366134 705798
rect 365514 691174 366134 705242
rect 365514 690618 365546 691174
rect 366102 690618 366134 691174
rect 365514 655174 366134 690618
rect 365514 654618 365546 655174
rect 366102 654618 366134 655174
rect 365514 619174 366134 654618
rect 365514 618618 365546 619174
rect 366102 618618 366134 619174
rect 365514 583174 366134 618618
rect 365514 582618 365546 583174
rect 366102 582618 366134 583174
rect 365514 547174 366134 582618
rect 365514 546618 365546 547174
rect 366102 546618 366134 547174
rect 365514 511174 366134 546618
rect 365514 510618 365546 511174
rect 366102 510618 366134 511174
rect 365514 475174 366134 510618
rect 365514 474618 365546 475174
rect 366102 474618 366134 475174
rect 365514 439174 366134 474618
rect 365514 438618 365546 439174
rect 366102 438618 366134 439174
rect 365514 403174 366134 438618
rect 365514 402618 365546 403174
rect 366102 402618 366134 403174
rect 365514 367174 366134 402618
rect 365514 366618 365546 367174
rect 366102 366618 366134 367174
rect 365514 331174 366134 366618
rect 369234 706758 369854 711590
rect 369234 706202 369266 706758
rect 369822 706202 369854 706758
rect 369234 694894 369854 706202
rect 369234 694338 369266 694894
rect 369822 694338 369854 694894
rect 369234 658894 369854 694338
rect 369234 658338 369266 658894
rect 369822 658338 369854 658894
rect 369234 622894 369854 658338
rect 369234 622338 369266 622894
rect 369822 622338 369854 622894
rect 369234 586894 369854 622338
rect 369234 586338 369266 586894
rect 369822 586338 369854 586894
rect 369234 550894 369854 586338
rect 369234 550338 369266 550894
rect 369822 550338 369854 550894
rect 369234 514894 369854 550338
rect 369234 514338 369266 514894
rect 369822 514338 369854 514894
rect 369234 478894 369854 514338
rect 369234 478338 369266 478894
rect 369822 478338 369854 478894
rect 369234 442894 369854 478338
rect 369234 442338 369266 442894
rect 369822 442338 369854 442894
rect 369234 406894 369854 442338
rect 369234 406338 369266 406894
rect 369822 406338 369854 406894
rect 369234 370894 369854 406338
rect 369234 370338 369266 370894
rect 369822 370338 369854 370894
rect 369234 354900 369854 370338
rect 372954 707718 373574 711590
rect 372954 707162 372986 707718
rect 373542 707162 373574 707718
rect 372954 698614 373574 707162
rect 372954 698058 372986 698614
rect 373542 698058 373574 698614
rect 372954 662614 373574 698058
rect 372954 662058 372986 662614
rect 373542 662058 373574 662614
rect 372954 626614 373574 662058
rect 372954 626058 372986 626614
rect 373542 626058 373574 626614
rect 372954 590614 373574 626058
rect 372954 590058 372986 590614
rect 373542 590058 373574 590614
rect 372954 554614 373574 590058
rect 372954 554058 372986 554614
rect 373542 554058 373574 554614
rect 372954 518614 373574 554058
rect 372954 518058 372986 518614
rect 373542 518058 373574 518614
rect 372954 482614 373574 518058
rect 372954 482058 372986 482614
rect 373542 482058 373574 482614
rect 372954 446614 373574 482058
rect 372954 446058 372986 446614
rect 373542 446058 373574 446614
rect 372954 410614 373574 446058
rect 372954 410058 372986 410614
rect 373542 410058 373574 410614
rect 372954 374614 373574 410058
rect 372954 374058 372986 374614
rect 373542 374058 373574 374614
rect 372954 338614 373574 374058
rect 372954 338058 372986 338614
rect 373542 338058 373574 338614
rect 365514 330618 365546 331174
rect 366102 330618 366134 331174
rect 365514 295174 366134 330618
rect 369488 331174 369808 331206
rect 369488 330938 369530 331174
rect 369766 330938 369808 331174
rect 369488 330854 369808 330938
rect 369488 330618 369530 330854
rect 369766 330618 369808 330854
rect 369488 330586 369808 330618
rect 372954 302614 373574 338058
rect 372954 302058 372986 302614
rect 373542 302058 373574 302614
rect 365514 294618 365546 295174
rect 366102 294618 366134 295174
rect 365514 259174 366134 294618
rect 369488 295174 369808 295206
rect 369488 294938 369530 295174
rect 369766 294938 369808 295174
rect 369488 294854 369808 294938
rect 369488 294618 369530 294854
rect 369766 294618 369808 294854
rect 369488 294586 369808 294618
rect 372954 266614 373574 302058
rect 372954 266058 372986 266614
rect 373542 266058 373574 266614
rect 365514 258618 365546 259174
rect 366102 258618 366134 259174
rect 365514 223174 366134 258618
rect 369488 259174 369808 259206
rect 369488 258938 369530 259174
rect 369766 258938 369808 259174
rect 369488 258854 369808 258938
rect 369488 258618 369530 258854
rect 369766 258618 369808 258854
rect 369488 258586 369808 258618
rect 372954 230614 373574 266058
rect 372954 230058 372986 230614
rect 373542 230058 373574 230614
rect 365514 222618 365546 223174
rect 366102 222618 366134 223174
rect 365514 187174 366134 222618
rect 369488 223174 369808 223206
rect 369488 222938 369530 223174
rect 369766 222938 369808 223174
rect 369488 222854 369808 222938
rect 369488 222618 369530 222854
rect 369766 222618 369808 222854
rect 369488 222586 369808 222618
rect 372954 194614 373574 230058
rect 372954 194058 372986 194614
rect 373542 194058 373574 194614
rect 365514 186618 365546 187174
rect 366102 186618 366134 187174
rect 365514 151174 366134 186618
rect 369488 187174 369808 187206
rect 369488 186938 369530 187174
rect 369766 186938 369808 187174
rect 369488 186854 369808 186938
rect 369488 186618 369530 186854
rect 369766 186618 369808 186854
rect 369488 186586 369808 186618
rect 372954 158614 373574 194058
rect 372954 158058 372986 158614
rect 373542 158058 373574 158614
rect 365514 150618 365546 151174
rect 366102 150618 366134 151174
rect 365514 115174 366134 150618
rect 369488 151174 369808 151206
rect 369488 150938 369530 151174
rect 369766 150938 369808 151174
rect 369488 150854 369808 150938
rect 369488 150618 369530 150854
rect 369766 150618 369808 150854
rect 369488 150586 369808 150618
rect 372954 122614 373574 158058
rect 372954 122058 372986 122614
rect 373542 122058 373574 122614
rect 365514 114618 365546 115174
rect 366102 114618 366134 115174
rect 365514 79174 366134 114618
rect 369488 115174 369808 115206
rect 369488 114938 369530 115174
rect 369766 114938 369808 115174
rect 369488 114854 369808 114938
rect 369488 114618 369530 114854
rect 369766 114618 369808 114854
rect 369488 114586 369808 114618
rect 372954 86614 373574 122058
rect 372954 86058 372986 86614
rect 373542 86058 373574 86614
rect 365514 78618 365546 79174
rect 366102 78618 366134 79174
rect 365514 43174 366134 78618
rect 369488 79174 369808 79206
rect 369488 78938 369530 79174
rect 369766 78938 369808 79174
rect 369488 78854 369808 78938
rect 369488 78618 369530 78854
rect 369766 78618 369808 78854
rect 369488 78586 369808 78618
rect 372954 50614 373574 86058
rect 372954 50058 372986 50614
rect 373542 50058 373574 50614
rect 365514 42618 365546 43174
rect 366102 42618 366134 43174
rect 365514 7174 366134 42618
rect 369488 43174 369808 43206
rect 369488 42938 369530 43174
rect 369766 42938 369808 43174
rect 369488 42854 369808 42938
rect 369488 42618 369530 42854
rect 369766 42618 369808 42854
rect 369488 42586 369808 42618
rect 372954 14614 373574 50058
rect 372954 14058 372986 14614
rect 373542 14058 373574 14614
rect 365514 6618 365546 7174
rect 366102 6618 366134 7174
rect 365514 -1306 366134 6618
rect 369488 7174 369808 7206
rect 369488 6938 369530 7174
rect 369766 6938 369808 7174
rect 369488 6854 369808 6938
rect 369488 6618 369530 6854
rect 369766 6618 369808 6854
rect 369488 6586 369808 6618
rect 365514 -1862 365546 -1306
rect 366102 -1862 366134 -1306
rect 365514 -7654 366134 -1862
rect 372954 -3226 373574 14058
rect 372954 -3782 372986 -3226
rect 373542 -3782 373574 -3226
rect 372954 -7654 373574 -3782
rect 376674 708678 377294 711590
rect 376674 708122 376706 708678
rect 377262 708122 377294 708678
rect 376674 666334 377294 708122
rect 376674 665778 376706 666334
rect 377262 665778 377294 666334
rect 376674 630334 377294 665778
rect 376674 629778 376706 630334
rect 377262 629778 377294 630334
rect 376674 594334 377294 629778
rect 376674 593778 376706 594334
rect 377262 593778 377294 594334
rect 376674 558334 377294 593778
rect 376674 557778 376706 558334
rect 377262 557778 377294 558334
rect 376674 522334 377294 557778
rect 376674 521778 376706 522334
rect 377262 521778 377294 522334
rect 376674 486334 377294 521778
rect 376674 485778 376706 486334
rect 377262 485778 377294 486334
rect 376674 450334 377294 485778
rect 376674 449778 376706 450334
rect 377262 449778 377294 450334
rect 376674 414334 377294 449778
rect 376674 413778 376706 414334
rect 377262 413778 377294 414334
rect 376674 378334 377294 413778
rect 376674 377778 376706 378334
rect 377262 377778 377294 378334
rect 376674 342334 377294 377778
rect 376674 341778 376706 342334
rect 377262 341778 377294 342334
rect 376674 306334 377294 341778
rect 376674 305778 376706 306334
rect 377262 305778 377294 306334
rect 376674 270334 377294 305778
rect 376674 269778 376706 270334
rect 377262 269778 377294 270334
rect 376674 234334 377294 269778
rect 376674 233778 376706 234334
rect 377262 233778 377294 234334
rect 376674 198334 377294 233778
rect 376674 197778 376706 198334
rect 377262 197778 377294 198334
rect 376674 162334 377294 197778
rect 376674 161778 376706 162334
rect 377262 161778 377294 162334
rect 376674 126334 377294 161778
rect 376674 125778 376706 126334
rect 377262 125778 377294 126334
rect 376674 90334 377294 125778
rect 376674 89778 376706 90334
rect 377262 89778 377294 90334
rect 376674 54334 377294 89778
rect 376674 53778 376706 54334
rect 377262 53778 377294 54334
rect 376674 18334 377294 53778
rect 376674 17778 376706 18334
rect 377262 17778 377294 18334
rect 376674 -4186 377294 17778
rect 376674 -4742 376706 -4186
rect 377262 -4742 377294 -4186
rect 376674 -7654 377294 -4742
rect 380394 709638 381014 711590
rect 380394 709082 380426 709638
rect 380982 709082 381014 709638
rect 380394 670054 381014 709082
rect 380394 669498 380426 670054
rect 380982 669498 381014 670054
rect 380394 634054 381014 669498
rect 380394 633498 380426 634054
rect 380982 633498 381014 634054
rect 380394 598054 381014 633498
rect 380394 597498 380426 598054
rect 380982 597498 381014 598054
rect 380394 562054 381014 597498
rect 380394 561498 380426 562054
rect 380982 561498 381014 562054
rect 380394 526054 381014 561498
rect 380394 525498 380426 526054
rect 380982 525498 381014 526054
rect 380394 490054 381014 525498
rect 380394 489498 380426 490054
rect 380982 489498 381014 490054
rect 380394 454054 381014 489498
rect 380394 453498 380426 454054
rect 380982 453498 381014 454054
rect 380394 418054 381014 453498
rect 380394 417498 380426 418054
rect 380982 417498 381014 418054
rect 380394 382054 381014 417498
rect 380394 381498 380426 382054
rect 380982 381498 381014 382054
rect 380394 346054 381014 381498
rect 380394 345498 380426 346054
rect 380982 345498 381014 346054
rect 380394 310054 381014 345498
rect 380394 309498 380426 310054
rect 380982 309498 381014 310054
rect 380394 274054 381014 309498
rect 380394 273498 380426 274054
rect 380982 273498 381014 274054
rect 380394 238054 381014 273498
rect 380394 237498 380426 238054
rect 380982 237498 381014 238054
rect 380394 202054 381014 237498
rect 380394 201498 380426 202054
rect 380982 201498 381014 202054
rect 380394 166054 381014 201498
rect 380394 165498 380426 166054
rect 380982 165498 381014 166054
rect 380394 130054 381014 165498
rect 380394 129498 380426 130054
rect 380982 129498 381014 130054
rect 380394 94054 381014 129498
rect 380394 93498 380426 94054
rect 380982 93498 381014 94054
rect 380394 58054 381014 93498
rect 380394 57498 380426 58054
rect 380982 57498 381014 58054
rect 380394 22054 381014 57498
rect 380394 21498 380426 22054
rect 380982 21498 381014 22054
rect 380394 -5146 381014 21498
rect 380394 -5702 380426 -5146
rect 380982 -5702 381014 -5146
rect 380394 -7654 381014 -5702
rect 384114 710598 384734 711590
rect 384114 710042 384146 710598
rect 384702 710042 384734 710598
rect 384114 673774 384734 710042
rect 384114 673218 384146 673774
rect 384702 673218 384734 673774
rect 384114 637774 384734 673218
rect 384114 637218 384146 637774
rect 384702 637218 384734 637774
rect 384114 601774 384734 637218
rect 384114 601218 384146 601774
rect 384702 601218 384734 601774
rect 384114 565774 384734 601218
rect 384114 565218 384146 565774
rect 384702 565218 384734 565774
rect 384114 529774 384734 565218
rect 384114 529218 384146 529774
rect 384702 529218 384734 529774
rect 384114 493774 384734 529218
rect 384114 493218 384146 493774
rect 384702 493218 384734 493774
rect 384114 457774 384734 493218
rect 384114 457218 384146 457774
rect 384702 457218 384734 457774
rect 384114 421774 384734 457218
rect 384114 421218 384146 421774
rect 384702 421218 384734 421774
rect 384114 385774 384734 421218
rect 384114 385218 384146 385774
rect 384702 385218 384734 385774
rect 384114 349774 384734 385218
rect 384114 349218 384146 349774
rect 384702 349218 384734 349774
rect 384114 313774 384734 349218
rect 387834 711558 388454 711590
rect 387834 711002 387866 711558
rect 388422 711002 388454 711558
rect 387834 677494 388454 711002
rect 387834 676938 387866 677494
rect 388422 676938 388454 677494
rect 387834 641494 388454 676938
rect 387834 640938 387866 641494
rect 388422 640938 388454 641494
rect 387834 605494 388454 640938
rect 387834 604938 387866 605494
rect 388422 604938 388454 605494
rect 387834 569494 388454 604938
rect 387834 568938 387866 569494
rect 388422 568938 388454 569494
rect 387834 533494 388454 568938
rect 387834 532938 387866 533494
rect 388422 532938 388454 533494
rect 387834 497494 388454 532938
rect 387834 496938 387866 497494
rect 388422 496938 388454 497494
rect 387834 461494 388454 496938
rect 387834 460938 387866 461494
rect 388422 460938 388454 461494
rect 387834 425494 388454 460938
rect 387834 424938 387866 425494
rect 388422 424938 388454 425494
rect 387834 389494 388454 424938
rect 387834 388938 387866 389494
rect 388422 388938 388454 389494
rect 387834 353494 388454 388938
rect 387834 352938 387866 353494
rect 388422 352938 388454 353494
rect 384848 327454 385168 327486
rect 384848 327218 384890 327454
rect 385126 327218 385168 327454
rect 384848 327134 385168 327218
rect 384848 326898 384890 327134
rect 385126 326898 385168 327134
rect 384848 326866 385168 326898
rect 384114 313218 384146 313774
rect 384702 313218 384734 313774
rect 384114 277774 384734 313218
rect 387834 317494 388454 352938
rect 387834 316938 387866 317494
rect 388422 316938 388454 317494
rect 384848 291454 385168 291486
rect 384848 291218 384890 291454
rect 385126 291218 385168 291454
rect 384848 291134 385168 291218
rect 384848 290898 384890 291134
rect 385126 290898 385168 291134
rect 384848 290866 385168 290898
rect 384114 277218 384146 277774
rect 384702 277218 384734 277774
rect 384114 241774 384734 277218
rect 387834 281494 388454 316938
rect 387834 280938 387866 281494
rect 388422 280938 388454 281494
rect 384848 255454 385168 255486
rect 384848 255218 384890 255454
rect 385126 255218 385168 255454
rect 384848 255134 385168 255218
rect 384848 254898 384890 255134
rect 385126 254898 385168 255134
rect 384848 254866 385168 254898
rect 384114 241218 384146 241774
rect 384702 241218 384734 241774
rect 384114 205774 384734 241218
rect 387834 245494 388454 280938
rect 387834 244938 387866 245494
rect 388422 244938 388454 245494
rect 384848 219454 385168 219486
rect 384848 219218 384890 219454
rect 385126 219218 385168 219454
rect 384848 219134 385168 219218
rect 384848 218898 384890 219134
rect 385126 218898 385168 219134
rect 384848 218866 385168 218898
rect 384114 205218 384146 205774
rect 384702 205218 384734 205774
rect 384114 169774 384734 205218
rect 387834 209494 388454 244938
rect 387834 208938 387866 209494
rect 388422 208938 388454 209494
rect 384848 183454 385168 183486
rect 384848 183218 384890 183454
rect 385126 183218 385168 183454
rect 384848 183134 385168 183218
rect 384848 182898 384890 183134
rect 385126 182898 385168 183134
rect 384848 182866 385168 182898
rect 384114 169218 384146 169774
rect 384702 169218 384734 169774
rect 384114 133774 384734 169218
rect 387834 173494 388454 208938
rect 387834 172938 387866 173494
rect 388422 172938 388454 173494
rect 384848 147454 385168 147486
rect 384848 147218 384890 147454
rect 385126 147218 385168 147454
rect 384848 147134 385168 147218
rect 384848 146898 384890 147134
rect 385126 146898 385168 147134
rect 384848 146866 385168 146898
rect 384114 133218 384146 133774
rect 384702 133218 384734 133774
rect 384114 97774 384734 133218
rect 387834 137494 388454 172938
rect 387834 136938 387866 137494
rect 388422 136938 388454 137494
rect 384848 111454 385168 111486
rect 384848 111218 384890 111454
rect 385126 111218 385168 111454
rect 384848 111134 385168 111218
rect 384848 110898 384890 111134
rect 385126 110898 385168 111134
rect 384848 110866 385168 110898
rect 384114 97218 384146 97774
rect 384702 97218 384734 97774
rect 384114 61774 384734 97218
rect 387834 101494 388454 136938
rect 387834 100938 387866 101494
rect 388422 100938 388454 101494
rect 384848 75454 385168 75486
rect 384848 75218 384890 75454
rect 385126 75218 385168 75454
rect 384848 75134 385168 75218
rect 384848 74898 384890 75134
rect 385126 74898 385168 75134
rect 384848 74866 385168 74898
rect 384114 61218 384146 61774
rect 384702 61218 384734 61774
rect 384114 25774 384734 61218
rect 387834 65494 388454 100938
rect 387834 64938 387866 65494
rect 388422 64938 388454 65494
rect 384848 39454 385168 39486
rect 384848 39218 384890 39454
rect 385126 39218 385168 39454
rect 384848 39134 385168 39218
rect 384848 38898 384890 39134
rect 385126 38898 385168 39134
rect 384848 38866 385168 38898
rect 384114 25218 384146 25774
rect 384702 25218 384734 25774
rect 384114 -6106 384734 25218
rect 384114 -6662 384146 -6106
rect 384702 -6662 384734 -6106
rect 384114 -7654 384734 -6662
rect 387834 29494 388454 64938
rect 387834 28938 387866 29494
rect 388422 28938 388454 29494
rect 387834 -7066 388454 28938
rect 387834 -7622 387866 -7066
rect 388422 -7622 388454 -7066
rect 387834 -7654 388454 -7622
rect 397794 704838 398414 711590
rect 397794 704282 397826 704838
rect 398382 704282 398414 704838
rect 397794 687454 398414 704282
rect 397794 686898 397826 687454
rect 398382 686898 398414 687454
rect 397794 651454 398414 686898
rect 397794 650898 397826 651454
rect 398382 650898 398414 651454
rect 397794 615454 398414 650898
rect 397794 614898 397826 615454
rect 398382 614898 398414 615454
rect 397794 579454 398414 614898
rect 397794 578898 397826 579454
rect 398382 578898 398414 579454
rect 397794 543454 398414 578898
rect 397794 542898 397826 543454
rect 398382 542898 398414 543454
rect 397794 507454 398414 542898
rect 397794 506898 397826 507454
rect 398382 506898 398414 507454
rect 397794 471454 398414 506898
rect 397794 470898 397826 471454
rect 398382 470898 398414 471454
rect 397794 435454 398414 470898
rect 397794 434898 397826 435454
rect 398382 434898 398414 435454
rect 397794 399454 398414 434898
rect 397794 398898 397826 399454
rect 398382 398898 398414 399454
rect 397794 363454 398414 398898
rect 397794 362898 397826 363454
rect 398382 362898 398414 363454
rect 397794 327454 398414 362898
rect 401514 705798 402134 711590
rect 401514 705242 401546 705798
rect 402102 705242 402134 705798
rect 401514 691174 402134 705242
rect 401514 690618 401546 691174
rect 402102 690618 402134 691174
rect 401514 655174 402134 690618
rect 401514 654618 401546 655174
rect 402102 654618 402134 655174
rect 401514 619174 402134 654618
rect 401514 618618 401546 619174
rect 402102 618618 402134 619174
rect 401514 583174 402134 618618
rect 401514 582618 401546 583174
rect 402102 582618 402134 583174
rect 401514 547174 402134 582618
rect 401514 546618 401546 547174
rect 402102 546618 402134 547174
rect 401514 511174 402134 546618
rect 401514 510618 401546 511174
rect 402102 510618 402134 511174
rect 401514 475174 402134 510618
rect 401514 474618 401546 475174
rect 402102 474618 402134 475174
rect 401514 439174 402134 474618
rect 401514 438618 401546 439174
rect 402102 438618 402134 439174
rect 401514 403174 402134 438618
rect 401514 402618 401546 403174
rect 402102 402618 402134 403174
rect 401514 367174 402134 402618
rect 401514 366618 401546 367174
rect 402102 366618 402134 367174
rect 400208 331174 400528 331206
rect 400208 330938 400250 331174
rect 400486 330938 400528 331174
rect 400208 330854 400528 330938
rect 400208 330618 400250 330854
rect 400486 330618 400528 330854
rect 400208 330586 400528 330618
rect 401514 331174 402134 366618
rect 401514 330618 401546 331174
rect 402102 330618 402134 331174
rect 397794 326898 397826 327454
rect 398382 326898 398414 327454
rect 397794 291454 398414 326898
rect 400208 295174 400528 295206
rect 400208 294938 400250 295174
rect 400486 294938 400528 295174
rect 400208 294854 400528 294938
rect 400208 294618 400250 294854
rect 400486 294618 400528 294854
rect 400208 294586 400528 294618
rect 401514 295174 402134 330618
rect 401514 294618 401546 295174
rect 402102 294618 402134 295174
rect 397794 290898 397826 291454
rect 398382 290898 398414 291454
rect 397794 255454 398414 290898
rect 400208 259174 400528 259206
rect 400208 258938 400250 259174
rect 400486 258938 400528 259174
rect 400208 258854 400528 258938
rect 400208 258618 400250 258854
rect 400486 258618 400528 258854
rect 400208 258586 400528 258618
rect 401514 259174 402134 294618
rect 401514 258618 401546 259174
rect 402102 258618 402134 259174
rect 397794 254898 397826 255454
rect 398382 254898 398414 255454
rect 397794 219454 398414 254898
rect 400208 223174 400528 223206
rect 400208 222938 400250 223174
rect 400486 222938 400528 223174
rect 400208 222854 400528 222938
rect 400208 222618 400250 222854
rect 400486 222618 400528 222854
rect 400208 222586 400528 222618
rect 401514 223174 402134 258618
rect 401514 222618 401546 223174
rect 402102 222618 402134 223174
rect 397794 218898 397826 219454
rect 398382 218898 398414 219454
rect 397794 183454 398414 218898
rect 400208 187174 400528 187206
rect 400208 186938 400250 187174
rect 400486 186938 400528 187174
rect 400208 186854 400528 186938
rect 400208 186618 400250 186854
rect 400486 186618 400528 186854
rect 400208 186586 400528 186618
rect 401514 187174 402134 222618
rect 401514 186618 401546 187174
rect 402102 186618 402134 187174
rect 397794 182898 397826 183454
rect 398382 182898 398414 183454
rect 397794 147454 398414 182898
rect 400208 151174 400528 151206
rect 400208 150938 400250 151174
rect 400486 150938 400528 151174
rect 400208 150854 400528 150938
rect 400208 150618 400250 150854
rect 400486 150618 400528 150854
rect 400208 150586 400528 150618
rect 401514 151174 402134 186618
rect 401514 150618 401546 151174
rect 402102 150618 402134 151174
rect 397794 146898 397826 147454
rect 398382 146898 398414 147454
rect 397794 111454 398414 146898
rect 400208 115174 400528 115206
rect 400208 114938 400250 115174
rect 400486 114938 400528 115174
rect 400208 114854 400528 114938
rect 400208 114618 400250 114854
rect 400486 114618 400528 114854
rect 400208 114586 400528 114618
rect 401514 115174 402134 150618
rect 401514 114618 401546 115174
rect 402102 114618 402134 115174
rect 397794 110898 397826 111454
rect 398382 110898 398414 111454
rect 397794 75454 398414 110898
rect 400208 79174 400528 79206
rect 400208 78938 400250 79174
rect 400486 78938 400528 79174
rect 400208 78854 400528 78938
rect 400208 78618 400250 78854
rect 400486 78618 400528 78854
rect 400208 78586 400528 78618
rect 401514 79174 402134 114618
rect 401514 78618 401546 79174
rect 402102 78618 402134 79174
rect 397794 74898 397826 75454
rect 398382 74898 398414 75454
rect 397794 39454 398414 74898
rect 400208 43174 400528 43206
rect 400208 42938 400250 43174
rect 400486 42938 400528 43174
rect 400208 42854 400528 42938
rect 400208 42618 400250 42854
rect 400486 42618 400528 42854
rect 400208 42586 400528 42618
rect 401514 43174 402134 78618
rect 401514 42618 401546 43174
rect 402102 42618 402134 43174
rect 397794 38898 397826 39454
rect 398382 38898 398414 39454
rect 397794 3454 398414 38898
rect 400208 7174 400528 7206
rect 400208 6938 400250 7174
rect 400486 6938 400528 7174
rect 400208 6854 400528 6938
rect 400208 6618 400250 6854
rect 400486 6618 400528 6854
rect 400208 6586 400528 6618
rect 401514 7174 402134 42618
rect 401514 6618 401546 7174
rect 402102 6618 402134 7174
rect 397794 2898 397826 3454
rect 398382 2898 398414 3454
rect 397794 -346 398414 2898
rect 397794 -902 397826 -346
rect 398382 -902 398414 -346
rect 397794 -7654 398414 -902
rect 401514 -1306 402134 6618
rect 401514 -1862 401546 -1306
rect 402102 -1862 402134 -1306
rect 401514 -7654 402134 -1862
rect 405234 706758 405854 711590
rect 405234 706202 405266 706758
rect 405822 706202 405854 706758
rect 405234 694894 405854 706202
rect 405234 694338 405266 694894
rect 405822 694338 405854 694894
rect 405234 658894 405854 694338
rect 405234 658338 405266 658894
rect 405822 658338 405854 658894
rect 405234 622894 405854 658338
rect 405234 622338 405266 622894
rect 405822 622338 405854 622894
rect 405234 586894 405854 622338
rect 405234 586338 405266 586894
rect 405822 586338 405854 586894
rect 405234 550894 405854 586338
rect 405234 550338 405266 550894
rect 405822 550338 405854 550894
rect 405234 514894 405854 550338
rect 405234 514338 405266 514894
rect 405822 514338 405854 514894
rect 405234 478894 405854 514338
rect 405234 478338 405266 478894
rect 405822 478338 405854 478894
rect 405234 442894 405854 478338
rect 405234 442338 405266 442894
rect 405822 442338 405854 442894
rect 405234 406894 405854 442338
rect 405234 406338 405266 406894
rect 405822 406338 405854 406894
rect 405234 370894 405854 406338
rect 405234 370338 405266 370894
rect 405822 370338 405854 370894
rect 405234 334894 405854 370338
rect 405234 334338 405266 334894
rect 405822 334338 405854 334894
rect 405234 298894 405854 334338
rect 405234 298338 405266 298894
rect 405822 298338 405854 298894
rect 405234 262894 405854 298338
rect 405234 262338 405266 262894
rect 405822 262338 405854 262894
rect 405234 226894 405854 262338
rect 405234 226338 405266 226894
rect 405822 226338 405854 226894
rect 405234 190894 405854 226338
rect 405234 190338 405266 190894
rect 405822 190338 405854 190894
rect 405234 154894 405854 190338
rect 405234 154338 405266 154894
rect 405822 154338 405854 154894
rect 405234 118894 405854 154338
rect 405234 118338 405266 118894
rect 405822 118338 405854 118894
rect 405234 82894 405854 118338
rect 405234 82338 405266 82894
rect 405822 82338 405854 82894
rect 405234 46894 405854 82338
rect 405234 46338 405266 46894
rect 405822 46338 405854 46894
rect 405234 10894 405854 46338
rect 405234 10338 405266 10894
rect 405822 10338 405854 10894
rect 405234 -2266 405854 10338
rect 405234 -2822 405266 -2266
rect 405822 -2822 405854 -2266
rect 405234 -7654 405854 -2822
rect 408954 707718 409574 711590
rect 408954 707162 408986 707718
rect 409542 707162 409574 707718
rect 408954 698614 409574 707162
rect 408954 698058 408986 698614
rect 409542 698058 409574 698614
rect 408954 662614 409574 698058
rect 408954 662058 408986 662614
rect 409542 662058 409574 662614
rect 408954 626614 409574 662058
rect 408954 626058 408986 626614
rect 409542 626058 409574 626614
rect 408954 590614 409574 626058
rect 408954 590058 408986 590614
rect 409542 590058 409574 590614
rect 408954 554614 409574 590058
rect 408954 554058 408986 554614
rect 409542 554058 409574 554614
rect 408954 518614 409574 554058
rect 408954 518058 408986 518614
rect 409542 518058 409574 518614
rect 408954 482614 409574 518058
rect 408954 482058 408986 482614
rect 409542 482058 409574 482614
rect 408954 446614 409574 482058
rect 408954 446058 408986 446614
rect 409542 446058 409574 446614
rect 408954 410614 409574 446058
rect 408954 410058 408986 410614
rect 409542 410058 409574 410614
rect 408954 374614 409574 410058
rect 408954 374058 408986 374614
rect 409542 374058 409574 374614
rect 408954 338614 409574 374058
rect 408954 338058 408986 338614
rect 409542 338058 409574 338614
rect 408954 302614 409574 338058
rect 408954 302058 408986 302614
rect 409542 302058 409574 302614
rect 408954 266614 409574 302058
rect 408954 266058 408986 266614
rect 409542 266058 409574 266614
rect 408954 230614 409574 266058
rect 408954 230058 408986 230614
rect 409542 230058 409574 230614
rect 408954 194614 409574 230058
rect 408954 194058 408986 194614
rect 409542 194058 409574 194614
rect 408954 158614 409574 194058
rect 408954 158058 408986 158614
rect 409542 158058 409574 158614
rect 408954 122614 409574 158058
rect 408954 122058 408986 122614
rect 409542 122058 409574 122614
rect 408954 86614 409574 122058
rect 408954 86058 408986 86614
rect 409542 86058 409574 86614
rect 408954 50614 409574 86058
rect 408954 50058 408986 50614
rect 409542 50058 409574 50614
rect 408954 14614 409574 50058
rect 408954 14058 408986 14614
rect 409542 14058 409574 14614
rect 408954 -3226 409574 14058
rect 408954 -3782 408986 -3226
rect 409542 -3782 409574 -3226
rect 408954 -7654 409574 -3782
rect 412674 708678 413294 711590
rect 412674 708122 412706 708678
rect 413262 708122 413294 708678
rect 412674 666334 413294 708122
rect 412674 665778 412706 666334
rect 413262 665778 413294 666334
rect 412674 630334 413294 665778
rect 412674 629778 412706 630334
rect 413262 629778 413294 630334
rect 412674 594334 413294 629778
rect 412674 593778 412706 594334
rect 413262 593778 413294 594334
rect 412674 558334 413294 593778
rect 412674 557778 412706 558334
rect 413262 557778 413294 558334
rect 412674 522334 413294 557778
rect 412674 521778 412706 522334
rect 413262 521778 413294 522334
rect 412674 486334 413294 521778
rect 412674 485778 412706 486334
rect 413262 485778 413294 486334
rect 412674 450334 413294 485778
rect 412674 449778 412706 450334
rect 413262 449778 413294 450334
rect 412674 414334 413294 449778
rect 412674 413778 412706 414334
rect 413262 413778 413294 414334
rect 412674 378334 413294 413778
rect 412674 377778 412706 378334
rect 413262 377778 413294 378334
rect 412674 342334 413294 377778
rect 412674 341778 412706 342334
rect 413262 341778 413294 342334
rect 412674 306334 413294 341778
rect 416394 709638 417014 711590
rect 416394 709082 416426 709638
rect 416982 709082 417014 709638
rect 416394 670054 417014 709082
rect 416394 669498 416426 670054
rect 416982 669498 417014 670054
rect 416394 634054 417014 669498
rect 416394 633498 416426 634054
rect 416982 633498 417014 634054
rect 416394 598054 417014 633498
rect 416394 597498 416426 598054
rect 416982 597498 417014 598054
rect 416394 562054 417014 597498
rect 416394 561498 416426 562054
rect 416982 561498 417014 562054
rect 416394 526054 417014 561498
rect 416394 525498 416426 526054
rect 416982 525498 417014 526054
rect 416394 490054 417014 525498
rect 416394 489498 416426 490054
rect 416982 489498 417014 490054
rect 416394 454054 417014 489498
rect 416394 453498 416426 454054
rect 416982 453498 417014 454054
rect 416394 418054 417014 453498
rect 416394 417498 416426 418054
rect 416982 417498 417014 418054
rect 416394 382054 417014 417498
rect 416394 381498 416426 382054
rect 416982 381498 417014 382054
rect 416394 346054 417014 381498
rect 416394 345498 416426 346054
rect 416982 345498 417014 346054
rect 415568 327454 415888 327486
rect 415568 327218 415610 327454
rect 415846 327218 415888 327454
rect 415568 327134 415888 327218
rect 415568 326898 415610 327134
rect 415846 326898 415888 327134
rect 415568 326866 415888 326898
rect 412674 305778 412706 306334
rect 413262 305778 413294 306334
rect 412674 270334 413294 305778
rect 416394 310054 417014 345498
rect 416394 309498 416426 310054
rect 416982 309498 417014 310054
rect 415568 291454 415888 291486
rect 415568 291218 415610 291454
rect 415846 291218 415888 291454
rect 415568 291134 415888 291218
rect 415568 290898 415610 291134
rect 415846 290898 415888 291134
rect 415568 290866 415888 290898
rect 412674 269778 412706 270334
rect 413262 269778 413294 270334
rect 412674 234334 413294 269778
rect 416394 274054 417014 309498
rect 416394 273498 416426 274054
rect 416982 273498 417014 274054
rect 415568 255454 415888 255486
rect 415568 255218 415610 255454
rect 415846 255218 415888 255454
rect 415568 255134 415888 255218
rect 415568 254898 415610 255134
rect 415846 254898 415888 255134
rect 415568 254866 415888 254898
rect 412674 233778 412706 234334
rect 413262 233778 413294 234334
rect 412674 198334 413294 233778
rect 416394 238054 417014 273498
rect 416394 237498 416426 238054
rect 416982 237498 417014 238054
rect 415568 219454 415888 219486
rect 415568 219218 415610 219454
rect 415846 219218 415888 219454
rect 415568 219134 415888 219218
rect 415568 218898 415610 219134
rect 415846 218898 415888 219134
rect 415568 218866 415888 218898
rect 412674 197778 412706 198334
rect 413262 197778 413294 198334
rect 412674 162334 413294 197778
rect 416394 202054 417014 237498
rect 416394 201498 416426 202054
rect 416982 201498 417014 202054
rect 415568 183454 415888 183486
rect 415568 183218 415610 183454
rect 415846 183218 415888 183454
rect 415568 183134 415888 183218
rect 415568 182898 415610 183134
rect 415846 182898 415888 183134
rect 415568 182866 415888 182898
rect 412674 161778 412706 162334
rect 413262 161778 413294 162334
rect 412674 126334 413294 161778
rect 416394 166054 417014 201498
rect 416394 165498 416426 166054
rect 416982 165498 417014 166054
rect 415568 147454 415888 147486
rect 415568 147218 415610 147454
rect 415846 147218 415888 147454
rect 415568 147134 415888 147218
rect 415568 146898 415610 147134
rect 415846 146898 415888 147134
rect 415568 146866 415888 146898
rect 412674 125778 412706 126334
rect 413262 125778 413294 126334
rect 412674 90334 413294 125778
rect 416394 130054 417014 165498
rect 416394 129498 416426 130054
rect 416982 129498 417014 130054
rect 415568 111454 415888 111486
rect 415568 111218 415610 111454
rect 415846 111218 415888 111454
rect 415568 111134 415888 111218
rect 415568 110898 415610 111134
rect 415846 110898 415888 111134
rect 415568 110866 415888 110898
rect 412674 89778 412706 90334
rect 413262 89778 413294 90334
rect 412674 54334 413294 89778
rect 416394 94054 417014 129498
rect 416394 93498 416426 94054
rect 416982 93498 417014 94054
rect 415568 75454 415888 75486
rect 415568 75218 415610 75454
rect 415846 75218 415888 75454
rect 415568 75134 415888 75218
rect 415568 74898 415610 75134
rect 415846 74898 415888 75134
rect 415568 74866 415888 74898
rect 412674 53778 412706 54334
rect 413262 53778 413294 54334
rect 412674 18334 413294 53778
rect 416394 58054 417014 93498
rect 416394 57498 416426 58054
rect 416982 57498 417014 58054
rect 415568 39454 415888 39486
rect 415568 39218 415610 39454
rect 415846 39218 415888 39454
rect 415568 39134 415888 39218
rect 415568 38898 415610 39134
rect 415846 38898 415888 39134
rect 415568 38866 415888 38898
rect 412674 17778 412706 18334
rect 413262 17778 413294 18334
rect 412674 -4186 413294 17778
rect 412674 -4742 412706 -4186
rect 413262 -4742 413294 -4186
rect 412674 -7654 413294 -4742
rect 416394 22054 417014 57498
rect 416394 21498 416426 22054
rect 416982 21498 417014 22054
rect 416394 -5146 417014 21498
rect 416394 -5702 416426 -5146
rect 416982 -5702 417014 -5146
rect 416394 -7654 417014 -5702
rect 420114 710598 420734 711590
rect 420114 710042 420146 710598
rect 420702 710042 420734 710598
rect 420114 673774 420734 710042
rect 420114 673218 420146 673774
rect 420702 673218 420734 673774
rect 420114 637774 420734 673218
rect 420114 637218 420146 637774
rect 420702 637218 420734 637774
rect 420114 601774 420734 637218
rect 420114 601218 420146 601774
rect 420702 601218 420734 601774
rect 420114 565774 420734 601218
rect 420114 565218 420146 565774
rect 420702 565218 420734 565774
rect 420114 529774 420734 565218
rect 420114 529218 420146 529774
rect 420702 529218 420734 529774
rect 420114 493774 420734 529218
rect 420114 493218 420146 493774
rect 420702 493218 420734 493774
rect 420114 457774 420734 493218
rect 420114 457218 420146 457774
rect 420702 457218 420734 457774
rect 420114 421774 420734 457218
rect 420114 421218 420146 421774
rect 420702 421218 420734 421774
rect 420114 385774 420734 421218
rect 420114 385218 420146 385774
rect 420702 385218 420734 385774
rect 420114 349774 420734 385218
rect 420114 349218 420146 349774
rect 420702 349218 420734 349774
rect 420114 313774 420734 349218
rect 420114 313218 420146 313774
rect 420702 313218 420734 313774
rect 420114 277774 420734 313218
rect 420114 277218 420146 277774
rect 420702 277218 420734 277774
rect 420114 241774 420734 277218
rect 420114 241218 420146 241774
rect 420702 241218 420734 241774
rect 420114 205774 420734 241218
rect 420114 205218 420146 205774
rect 420702 205218 420734 205774
rect 420114 169774 420734 205218
rect 420114 169218 420146 169774
rect 420702 169218 420734 169774
rect 420114 133774 420734 169218
rect 420114 133218 420146 133774
rect 420702 133218 420734 133774
rect 420114 97774 420734 133218
rect 420114 97218 420146 97774
rect 420702 97218 420734 97774
rect 420114 61774 420734 97218
rect 420114 61218 420146 61774
rect 420702 61218 420734 61774
rect 420114 25774 420734 61218
rect 420114 25218 420146 25774
rect 420702 25218 420734 25774
rect 420114 -6106 420734 25218
rect 420114 -6662 420146 -6106
rect 420702 -6662 420734 -6106
rect 420114 -7654 420734 -6662
rect 423834 711558 424454 711590
rect 423834 711002 423866 711558
rect 424422 711002 424454 711558
rect 423834 677494 424454 711002
rect 423834 676938 423866 677494
rect 424422 676938 424454 677494
rect 423834 641494 424454 676938
rect 423834 640938 423866 641494
rect 424422 640938 424454 641494
rect 423834 605494 424454 640938
rect 423834 604938 423866 605494
rect 424422 604938 424454 605494
rect 423834 569494 424454 604938
rect 423834 568938 423866 569494
rect 424422 568938 424454 569494
rect 423834 533494 424454 568938
rect 423834 532938 423866 533494
rect 424422 532938 424454 533494
rect 423834 497494 424454 532938
rect 423834 496938 423866 497494
rect 424422 496938 424454 497494
rect 423834 461494 424454 496938
rect 423834 460938 423866 461494
rect 424422 460938 424454 461494
rect 423834 425494 424454 460938
rect 423834 424938 423866 425494
rect 424422 424938 424454 425494
rect 423834 389494 424454 424938
rect 423834 388938 423866 389494
rect 424422 388938 424454 389494
rect 423834 353494 424454 388938
rect 423834 352938 423866 353494
rect 424422 352938 424454 353494
rect 423834 317494 424454 352938
rect 433794 704838 434414 711590
rect 433794 704282 433826 704838
rect 434382 704282 434414 704838
rect 433794 687454 434414 704282
rect 433794 686898 433826 687454
rect 434382 686898 434414 687454
rect 433794 651454 434414 686898
rect 433794 650898 433826 651454
rect 434382 650898 434414 651454
rect 433794 615454 434414 650898
rect 433794 614898 433826 615454
rect 434382 614898 434414 615454
rect 433794 579454 434414 614898
rect 433794 578898 433826 579454
rect 434382 578898 434414 579454
rect 433794 543454 434414 578898
rect 433794 542898 433826 543454
rect 434382 542898 434414 543454
rect 433794 507454 434414 542898
rect 433794 506898 433826 507454
rect 434382 506898 434414 507454
rect 433794 471454 434414 506898
rect 433794 470898 433826 471454
rect 434382 470898 434414 471454
rect 433794 435454 434414 470898
rect 433794 434898 433826 435454
rect 434382 434898 434414 435454
rect 433794 399454 434414 434898
rect 433794 398898 433826 399454
rect 434382 398898 434414 399454
rect 433794 363454 434414 398898
rect 433794 362898 433826 363454
rect 434382 362898 434414 363454
rect 430928 331174 431248 331206
rect 430928 330938 430970 331174
rect 431206 330938 431248 331174
rect 430928 330854 431248 330938
rect 430928 330618 430970 330854
rect 431206 330618 431248 330854
rect 430928 330586 431248 330618
rect 423834 316938 423866 317494
rect 424422 316938 424454 317494
rect 423834 281494 424454 316938
rect 433794 327454 434414 362898
rect 433794 326898 433826 327454
rect 434382 326898 434414 327454
rect 430928 295174 431248 295206
rect 430928 294938 430970 295174
rect 431206 294938 431248 295174
rect 430928 294854 431248 294938
rect 430928 294618 430970 294854
rect 431206 294618 431248 294854
rect 430928 294586 431248 294618
rect 423834 280938 423866 281494
rect 424422 280938 424454 281494
rect 423834 245494 424454 280938
rect 433794 291454 434414 326898
rect 433794 290898 433826 291454
rect 434382 290898 434414 291454
rect 430928 259174 431248 259206
rect 430928 258938 430970 259174
rect 431206 258938 431248 259174
rect 430928 258854 431248 258938
rect 430928 258618 430970 258854
rect 431206 258618 431248 258854
rect 430928 258586 431248 258618
rect 423834 244938 423866 245494
rect 424422 244938 424454 245494
rect 423834 209494 424454 244938
rect 433794 255454 434414 290898
rect 433794 254898 433826 255454
rect 434382 254898 434414 255454
rect 430928 223174 431248 223206
rect 430928 222938 430970 223174
rect 431206 222938 431248 223174
rect 430928 222854 431248 222938
rect 430928 222618 430970 222854
rect 431206 222618 431248 222854
rect 430928 222586 431248 222618
rect 423834 208938 423866 209494
rect 424422 208938 424454 209494
rect 423834 173494 424454 208938
rect 433794 219454 434414 254898
rect 433794 218898 433826 219454
rect 434382 218898 434414 219454
rect 430928 187174 431248 187206
rect 430928 186938 430970 187174
rect 431206 186938 431248 187174
rect 430928 186854 431248 186938
rect 430928 186618 430970 186854
rect 431206 186618 431248 186854
rect 430928 186586 431248 186618
rect 423834 172938 423866 173494
rect 424422 172938 424454 173494
rect 423834 137494 424454 172938
rect 433794 183454 434414 218898
rect 433794 182898 433826 183454
rect 434382 182898 434414 183454
rect 430928 151174 431248 151206
rect 430928 150938 430970 151174
rect 431206 150938 431248 151174
rect 430928 150854 431248 150938
rect 430928 150618 430970 150854
rect 431206 150618 431248 150854
rect 430928 150586 431248 150618
rect 423834 136938 423866 137494
rect 424422 136938 424454 137494
rect 423834 101494 424454 136938
rect 433794 147454 434414 182898
rect 433794 146898 433826 147454
rect 434382 146898 434414 147454
rect 430928 115174 431248 115206
rect 430928 114938 430970 115174
rect 431206 114938 431248 115174
rect 430928 114854 431248 114938
rect 430928 114618 430970 114854
rect 431206 114618 431248 114854
rect 430928 114586 431248 114618
rect 423834 100938 423866 101494
rect 424422 100938 424454 101494
rect 423834 65494 424454 100938
rect 433794 111454 434414 146898
rect 433794 110898 433826 111454
rect 434382 110898 434414 111454
rect 430928 79174 431248 79206
rect 430928 78938 430970 79174
rect 431206 78938 431248 79174
rect 430928 78854 431248 78938
rect 430928 78618 430970 78854
rect 431206 78618 431248 78854
rect 430928 78586 431248 78618
rect 423834 64938 423866 65494
rect 424422 64938 424454 65494
rect 423834 29494 424454 64938
rect 433794 75454 434414 110898
rect 433794 74898 433826 75454
rect 434382 74898 434414 75454
rect 430928 43174 431248 43206
rect 430928 42938 430970 43174
rect 431206 42938 431248 43174
rect 430928 42854 431248 42938
rect 430928 42618 430970 42854
rect 431206 42618 431248 42854
rect 430928 42586 431248 42618
rect 423834 28938 423866 29494
rect 424422 28938 424454 29494
rect 423834 -7066 424454 28938
rect 433794 39454 434414 74898
rect 433794 38898 433826 39454
rect 434382 38898 434414 39454
rect 430928 7174 431248 7206
rect 430928 6938 430970 7174
rect 431206 6938 431248 7174
rect 430928 6854 431248 6938
rect 430928 6618 430970 6854
rect 431206 6618 431248 6854
rect 430928 6586 431248 6618
rect 423834 -7622 423866 -7066
rect 424422 -7622 424454 -7066
rect 423834 -7654 424454 -7622
rect 433794 3454 434414 38898
rect 433794 2898 433826 3454
rect 434382 2898 434414 3454
rect 433794 -346 434414 2898
rect 433794 -902 433826 -346
rect 434382 -902 434414 -346
rect 433794 -7654 434414 -902
rect 437514 705798 438134 711590
rect 437514 705242 437546 705798
rect 438102 705242 438134 705798
rect 437514 691174 438134 705242
rect 437514 690618 437546 691174
rect 438102 690618 438134 691174
rect 437514 655174 438134 690618
rect 437514 654618 437546 655174
rect 438102 654618 438134 655174
rect 437514 619174 438134 654618
rect 437514 618618 437546 619174
rect 438102 618618 438134 619174
rect 437514 583174 438134 618618
rect 437514 582618 437546 583174
rect 438102 582618 438134 583174
rect 437514 547174 438134 582618
rect 437514 546618 437546 547174
rect 438102 546618 438134 547174
rect 437514 511174 438134 546618
rect 437514 510618 437546 511174
rect 438102 510618 438134 511174
rect 437514 475174 438134 510618
rect 437514 474618 437546 475174
rect 438102 474618 438134 475174
rect 437514 439174 438134 474618
rect 437514 438618 437546 439174
rect 438102 438618 438134 439174
rect 437514 403174 438134 438618
rect 437514 402618 437546 403174
rect 438102 402618 438134 403174
rect 437514 367174 438134 402618
rect 437514 366618 437546 367174
rect 438102 366618 438134 367174
rect 437514 331174 438134 366618
rect 437514 330618 437546 331174
rect 438102 330618 438134 331174
rect 437514 295174 438134 330618
rect 437514 294618 437546 295174
rect 438102 294618 438134 295174
rect 437514 259174 438134 294618
rect 437514 258618 437546 259174
rect 438102 258618 438134 259174
rect 437514 223174 438134 258618
rect 437514 222618 437546 223174
rect 438102 222618 438134 223174
rect 437514 187174 438134 222618
rect 437514 186618 437546 187174
rect 438102 186618 438134 187174
rect 437514 151174 438134 186618
rect 437514 150618 437546 151174
rect 438102 150618 438134 151174
rect 437514 115174 438134 150618
rect 437514 114618 437546 115174
rect 438102 114618 438134 115174
rect 437514 79174 438134 114618
rect 437514 78618 437546 79174
rect 438102 78618 438134 79174
rect 437514 43174 438134 78618
rect 437514 42618 437546 43174
rect 438102 42618 438134 43174
rect 437514 7174 438134 42618
rect 437514 6618 437546 7174
rect 438102 6618 438134 7174
rect 437514 -1306 438134 6618
rect 437514 -1862 437546 -1306
rect 438102 -1862 438134 -1306
rect 437514 -7654 438134 -1862
rect 441234 706758 441854 711590
rect 441234 706202 441266 706758
rect 441822 706202 441854 706758
rect 441234 694894 441854 706202
rect 441234 694338 441266 694894
rect 441822 694338 441854 694894
rect 441234 658894 441854 694338
rect 441234 658338 441266 658894
rect 441822 658338 441854 658894
rect 441234 622894 441854 658338
rect 441234 622338 441266 622894
rect 441822 622338 441854 622894
rect 441234 586894 441854 622338
rect 441234 586338 441266 586894
rect 441822 586338 441854 586894
rect 441234 550894 441854 586338
rect 441234 550338 441266 550894
rect 441822 550338 441854 550894
rect 441234 514894 441854 550338
rect 441234 514338 441266 514894
rect 441822 514338 441854 514894
rect 441234 478894 441854 514338
rect 441234 478338 441266 478894
rect 441822 478338 441854 478894
rect 441234 442894 441854 478338
rect 441234 442338 441266 442894
rect 441822 442338 441854 442894
rect 441234 406894 441854 442338
rect 441234 406338 441266 406894
rect 441822 406338 441854 406894
rect 441234 370894 441854 406338
rect 441234 370338 441266 370894
rect 441822 370338 441854 370894
rect 441234 334894 441854 370338
rect 441234 334338 441266 334894
rect 441822 334338 441854 334894
rect 441234 298894 441854 334338
rect 441234 298338 441266 298894
rect 441822 298338 441854 298894
rect 441234 262894 441854 298338
rect 441234 262338 441266 262894
rect 441822 262338 441854 262894
rect 441234 226894 441854 262338
rect 441234 226338 441266 226894
rect 441822 226338 441854 226894
rect 441234 190894 441854 226338
rect 441234 190338 441266 190894
rect 441822 190338 441854 190894
rect 441234 154894 441854 190338
rect 441234 154338 441266 154894
rect 441822 154338 441854 154894
rect 441234 118894 441854 154338
rect 441234 118338 441266 118894
rect 441822 118338 441854 118894
rect 441234 82894 441854 118338
rect 441234 82338 441266 82894
rect 441822 82338 441854 82894
rect 441234 46894 441854 82338
rect 441234 46338 441266 46894
rect 441822 46338 441854 46894
rect 441234 10894 441854 46338
rect 441234 10338 441266 10894
rect 441822 10338 441854 10894
rect 441234 -2266 441854 10338
rect 441234 -2822 441266 -2266
rect 441822 -2822 441854 -2266
rect 441234 -7654 441854 -2822
rect 444954 707718 445574 711590
rect 444954 707162 444986 707718
rect 445542 707162 445574 707718
rect 444954 698614 445574 707162
rect 444954 698058 444986 698614
rect 445542 698058 445574 698614
rect 444954 662614 445574 698058
rect 444954 662058 444986 662614
rect 445542 662058 445574 662614
rect 444954 626614 445574 662058
rect 444954 626058 444986 626614
rect 445542 626058 445574 626614
rect 444954 590614 445574 626058
rect 444954 590058 444986 590614
rect 445542 590058 445574 590614
rect 444954 554614 445574 590058
rect 444954 554058 444986 554614
rect 445542 554058 445574 554614
rect 444954 518614 445574 554058
rect 444954 518058 444986 518614
rect 445542 518058 445574 518614
rect 444954 482614 445574 518058
rect 444954 482058 444986 482614
rect 445542 482058 445574 482614
rect 444954 446614 445574 482058
rect 444954 446058 444986 446614
rect 445542 446058 445574 446614
rect 444954 410614 445574 446058
rect 444954 410058 444986 410614
rect 445542 410058 445574 410614
rect 444954 374614 445574 410058
rect 444954 374058 444986 374614
rect 445542 374058 445574 374614
rect 444954 338614 445574 374058
rect 444954 338058 444986 338614
rect 445542 338058 445574 338614
rect 444954 302614 445574 338058
rect 448674 708678 449294 711590
rect 448674 708122 448706 708678
rect 449262 708122 449294 708678
rect 448674 666334 449294 708122
rect 448674 665778 448706 666334
rect 449262 665778 449294 666334
rect 448674 630334 449294 665778
rect 448674 629778 448706 630334
rect 449262 629778 449294 630334
rect 448674 594334 449294 629778
rect 448674 593778 448706 594334
rect 449262 593778 449294 594334
rect 448674 558334 449294 593778
rect 448674 557778 448706 558334
rect 449262 557778 449294 558334
rect 448674 522334 449294 557778
rect 448674 521778 448706 522334
rect 449262 521778 449294 522334
rect 448674 486334 449294 521778
rect 448674 485778 448706 486334
rect 449262 485778 449294 486334
rect 448674 450334 449294 485778
rect 448674 449778 448706 450334
rect 449262 449778 449294 450334
rect 448674 414334 449294 449778
rect 448674 413778 448706 414334
rect 449262 413778 449294 414334
rect 448674 378334 449294 413778
rect 448674 377778 448706 378334
rect 449262 377778 449294 378334
rect 448674 342334 449294 377778
rect 448674 341778 448706 342334
rect 449262 341778 449294 342334
rect 446288 327454 446608 327486
rect 446288 327218 446330 327454
rect 446566 327218 446608 327454
rect 446288 327134 446608 327218
rect 446288 326898 446330 327134
rect 446566 326898 446608 327134
rect 446288 326866 446608 326898
rect 444954 302058 444986 302614
rect 445542 302058 445574 302614
rect 444954 266614 445574 302058
rect 448674 306334 449294 341778
rect 448674 305778 448706 306334
rect 449262 305778 449294 306334
rect 446288 291454 446608 291486
rect 446288 291218 446330 291454
rect 446566 291218 446608 291454
rect 446288 291134 446608 291218
rect 446288 290898 446330 291134
rect 446566 290898 446608 291134
rect 446288 290866 446608 290898
rect 444954 266058 444986 266614
rect 445542 266058 445574 266614
rect 444954 230614 445574 266058
rect 448674 270334 449294 305778
rect 448674 269778 448706 270334
rect 449262 269778 449294 270334
rect 446288 255454 446608 255486
rect 446288 255218 446330 255454
rect 446566 255218 446608 255454
rect 446288 255134 446608 255218
rect 446288 254898 446330 255134
rect 446566 254898 446608 255134
rect 446288 254866 446608 254898
rect 444954 230058 444986 230614
rect 445542 230058 445574 230614
rect 444954 194614 445574 230058
rect 448674 234334 449294 269778
rect 448674 233778 448706 234334
rect 449262 233778 449294 234334
rect 446288 219454 446608 219486
rect 446288 219218 446330 219454
rect 446566 219218 446608 219454
rect 446288 219134 446608 219218
rect 446288 218898 446330 219134
rect 446566 218898 446608 219134
rect 446288 218866 446608 218898
rect 444954 194058 444986 194614
rect 445542 194058 445574 194614
rect 444954 158614 445574 194058
rect 448674 198334 449294 233778
rect 448674 197778 448706 198334
rect 449262 197778 449294 198334
rect 446288 183454 446608 183486
rect 446288 183218 446330 183454
rect 446566 183218 446608 183454
rect 446288 183134 446608 183218
rect 446288 182898 446330 183134
rect 446566 182898 446608 183134
rect 446288 182866 446608 182898
rect 444954 158058 444986 158614
rect 445542 158058 445574 158614
rect 444954 122614 445574 158058
rect 448674 162334 449294 197778
rect 448674 161778 448706 162334
rect 449262 161778 449294 162334
rect 446288 147454 446608 147486
rect 446288 147218 446330 147454
rect 446566 147218 446608 147454
rect 446288 147134 446608 147218
rect 446288 146898 446330 147134
rect 446566 146898 446608 147134
rect 446288 146866 446608 146898
rect 444954 122058 444986 122614
rect 445542 122058 445574 122614
rect 444954 86614 445574 122058
rect 448674 126334 449294 161778
rect 448674 125778 448706 126334
rect 449262 125778 449294 126334
rect 446288 111454 446608 111486
rect 446288 111218 446330 111454
rect 446566 111218 446608 111454
rect 446288 111134 446608 111218
rect 446288 110898 446330 111134
rect 446566 110898 446608 111134
rect 446288 110866 446608 110898
rect 444954 86058 444986 86614
rect 445542 86058 445574 86614
rect 444954 50614 445574 86058
rect 448674 90334 449294 125778
rect 448674 89778 448706 90334
rect 449262 89778 449294 90334
rect 446288 75454 446608 75486
rect 446288 75218 446330 75454
rect 446566 75218 446608 75454
rect 446288 75134 446608 75218
rect 446288 74898 446330 75134
rect 446566 74898 446608 75134
rect 446288 74866 446608 74898
rect 444954 50058 444986 50614
rect 445542 50058 445574 50614
rect 444954 14614 445574 50058
rect 448674 54334 449294 89778
rect 448674 53778 448706 54334
rect 449262 53778 449294 54334
rect 446288 39454 446608 39486
rect 446288 39218 446330 39454
rect 446566 39218 446608 39454
rect 446288 39134 446608 39218
rect 446288 38898 446330 39134
rect 446566 38898 446608 39134
rect 446288 38866 446608 38898
rect 444954 14058 444986 14614
rect 445542 14058 445574 14614
rect 444954 -3226 445574 14058
rect 444954 -3782 444986 -3226
rect 445542 -3782 445574 -3226
rect 444954 -7654 445574 -3782
rect 448674 18334 449294 53778
rect 448674 17778 448706 18334
rect 449262 17778 449294 18334
rect 448674 -4186 449294 17778
rect 448674 -4742 448706 -4186
rect 449262 -4742 449294 -4186
rect 448674 -7654 449294 -4742
rect 452394 709638 453014 711590
rect 452394 709082 452426 709638
rect 452982 709082 453014 709638
rect 452394 670054 453014 709082
rect 452394 669498 452426 670054
rect 452982 669498 453014 670054
rect 452394 634054 453014 669498
rect 452394 633498 452426 634054
rect 452982 633498 453014 634054
rect 452394 598054 453014 633498
rect 452394 597498 452426 598054
rect 452982 597498 453014 598054
rect 452394 562054 453014 597498
rect 452394 561498 452426 562054
rect 452982 561498 453014 562054
rect 452394 526054 453014 561498
rect 452394 525498 452426 526054
rect 452982 525498 453014 526054
rect 452394 490054 453014 525498
rect 452394 489498 452426 490054
rect 452982 489498 453014 490054
rect 452394 454054 453014 489498
rect 452394 453498 452426 454054
rect 452982 453498 453014 454054
rect 452394 418054 453014 453498
rect 452394 417498 452426 418054
rect 452982 417498 453014 418054
rect 452394 382054 453014 417498
rect 452394 381498 452426 382054
rect 452982 381498 453014 382054
rect 452394 346054 453014 381498
rect 452394 345498 452426 346054
rect 452982 345498 453014 346054
rect 452394 310054 453014 345498
rect 452394 309498 452426 310054
rect 452982 309498 453014 310054
rect 452394 274054 453014 309498
rect 452394 273498 452426 274054
rect 452982 273498 453014 274054
rect 452394 238054 453014 273498
rect 452394 237498 452426 238054
rect 452982 237498 453014 238054
rect 452394 202054 453014 237498
rect 452394 201498 452426 202054
rect 452982 201498 453014 202054
rect 452394 166054 453014 201498
rect 452394 165498 452426 166054
rect 452982 165498 453014 166054
rect 452394 130054 453014 165498
rect 452394 129498 452426 130054
rect 452982 129498 453014 130054
rect 452394 94054 453014 129498
rect 452394 93498 452426 94054
rect 452982 93498 453014 94054
rect 452394 58054 453014 93498
rect 452394 57498 452426 58054
rect 452982 57498 453014 58054
rect 452394 22054 453014 57498
rect 452394 21498 452426 22054
rect 452982 21498 453014 22054
rect 452394 -5146 453014 21498
rect 452394 -5702 452426 -5146
rect 452982 -5702 453014 -5146
rect 452394 -7654 453014 -5702
rect 456114 710598 456734 711590
rect 456114 710042 456146 710598
rect 456702 710042 456734 710598
rect 456114 673774 456734 710042
rect 456114 673218 456146 673774
rect 456702 673218 456734 673774
rect 456114 637774 456734 673218
rect 456114 637218 456146 637774
rect 456702 637218 456734 637774
rect 456114 601774 456734 637218
rect 456114 601218 456146 601774
rect 456702 601218 456734 601774
rect 456114 565774 456734 601218
rect 456114 565218 456146 565774
rect 456702 565218 456734 565774
rect 456114 529774 456734 565218
rect 456114 529218 456146 529774
rect 456702 529218 456734 529774
rect 456114 493774 456734 529218
rect 456114 493218 456146 493774
rect 456702 493218 456734 493774
rect 456114 457774 456734 493218
rect 456114 457218 456146 457774
rect 456702 457218 456734 457774
rect 456114 421774 456734 457218
rect 456114 421218 456146 421774
rect 456702 421218 456734 421774
rect 456114 385774 456734 421218
rect 456114 385218 456146 385774
rect 456702 385218 456734 385774
rect 456114 349774 456734 385218
rect 456114 349218 456146 349774
rect 456702 349218 456734 349774
rect 456114 313774 456734 349218
rect 456114 313218 456146 313774
rect 456702 313218 456734 313774
rect 456114 277774 456734 313218
rect 456114 277218 456146 277774
rect 456702 277218 456734 277774
rect 456114 241774 456734 277218
rect 456114 241218 456146 241774
rect 456702 241218 456734 241774
rect 456114 205774 456734 241218
rect 456114 205218 456146 205774
rect 456702 205218 456734 205774
rect 456114 169774 456734 205218
rect 456114 169218 456146 169774
rect 456702 169218 456734 169774
rect 456114 133774 456734 169218
rect 456114 133218 456146 133774
rect 456702 133218 456734 133774
rect 456114 97774 456734 133218
rect 456114 97218 456146 97774
rect 456702 97218 456734 97774
rect 456114 61774 456734 97218
rect 456114 61218 456146 61774
rect 456702 61218 456734 61774
rect 456114 25774 456734 61218
rect 456114 25218 456146 25774
rect 456702 25218 456734 25774
rect 456114 -6106 456734 25218
rect 456114 -6662 456146 -6106
rect 456702 -6662 456734 -6106
rect 456114 -7654 456734 -6662
rect 459834 711558 460454 711590
rect 459834 711002 459866 711558
rect 460422 711002 460454 711558
rect 459834 677494 460454 711002
rect 459834 676938 459866 677494
rect 460422 676938 460454 677494
rect 459834 641494 460454 676938
rect 459834 640938 459866 641494
rect 460422 640938 460454 641494
rect 459834 605494 460454 640938
rect 459834 604938 459866 605494
rect 460422 604938 460454 605494
rect 459834 569494 460454 604938
rect 459834 568938 459866 569494
rect 460422 568938 460454 569494
rect 459834 533494 460454 568938
rect 459834 532938 459866 533494
rect 460422 532938 460454 533494
rect 459834 497494 460454 532938
rect 459834 496938 459866 497494
rect 460422 496938 460454 497494
rect 459834 461494 460454 496938
rect 459834 460938 459866 461494
rect 460422 460938 460454 461494
rect 459834 425494 460454 460938
rect 459834 424938 459866 425494
rect 460422 424938 460454 425494
rect 459834 389494 460454 424938
rect 459834 388938 459866 389494
rect 460422 388938 460454 389494
rect 459834 353494 460454 388938
rect 459834 352938 459866 353494
rect 460422 352938 460454 353494
rect 459834 317494 460454 352938
rect 469794 704838 470414 711590
rect 469794 704282 469826 704838
rect 470382 704282 470414 704838
rect 469794 687454 470414 704282
rect 469794 686898 469826 687454
rect 470382 686898 470414 687454
rect 469794 651454 470414 686898
rect 469794 650898 469826 651454
rect 470382 650898 470414 651454
rect 469794 615454 470414 650898
rect 469794 614898 469826 615454
rect 470382 614898 470414 615454
rect 469794 579454 470414 614898
rect 469794 578898 469826 579454
rect 470382 578898 470414 579454
rect 469794 543454 470414 578898
rect 469794 542898 469826 543454
rect 470382 542898 470414 543454
rect 469794 507454 470414 542898
rect 469794 506898 469826 507454
rect 470382 506898 470414 507454
rect 469794 471454 470414 506898
rect 469794 470898 469826 471454
rect 470382 470898 470414 471454
rect 469794 435454 470414 470898
rect 469794 434898 469826 435454
rect 470382 434898 470414 435454
rect 469794 399454 470414 434898
rect 469794 398898 469826 399454
rect 470382 398898 470414 399454
rect 469794 363454 470414 398898
rect 469794 362898 469826 363454
rect 470382 362898 470414 363454
rect 461648 331174 461968 331206
rect 461648 330938 461690 331174
rect 461926 330938 461968 331174
rect 461648 330854 461968 330938
rect 461648 330618 461690 330854
rect 461926 330618 461968 330854
rect 461648 330586 461968 330618
rect 459834 316938 459866 317494
rect 460422 316938 460454 317494
rect 459834 281494 460454 316938
rect 469794 327454 470414 362898
rect 469794 326898 469826 327454
rect 470382 326898 470414 327454
rect 461648 295174 461968 295206
rect 461648 294938 461690 295174
rect 461926 294938 461968 295174
rect 461648 294854 461968 294938
rect 461648 294618 461690 294854
rect 461926 294618 461968 294854
rect 461648 294586 461968 294618
rect 459834 280938 459866 281494
rect 460422 280938 460454 281494
rect 459834 245494 460454 280938
rect 469794 291454 470414 326898
rect 469794 290898 469826 291454
rect 470382 290898 470414 291454
rect 461648 259174 461968 259206
rect 461648 258938 461690 259174
rect 461926 258938 461968 259174
rect 461648 258854 461968 258938
rect 461648 258618 461690 258854
rect 461926 258618 461968 258854
rect 461648 258586 461968 258618
rect 459834 244938 459866 245494
rect 460422 244938 460454 245494
rect 459834 209494 460454 244938
rect 469794 255454 470414 290898
rect 469794 254898 469826 255454
rect 470382 254898 470414 255454
rect 461648 223174 461968 223206
rect 461648 222938 461690 223174
rect 461926 222938 461968 223174
rect 461648 222854 461968 222938
rect 461648 222618 461690 222854
rect 461926 222618 461968 222854
rect 461648 222586 461968 222618
rect 459834 208938 459866 209494
rect 460422 208938 460454 209494
rect 459834 173494 460454 208938
rect 469794 219454 470414 254898
rect 469794 218898 469826 219454
rect 470382 218898 470414 219454
rect 461648 187174 461968 187206
rect 461648 186938 461690 187174
rect 461926 186938 461968 187174
rect 461648 186854 461968 186938
rect 461648 186618 461690 186854
rect 461926 186618 461968 186854
rect 461648 186586 461968 186618
rect 459834 172938 459866 173494
rect 460422 172938 460454 173494
rect 459834 137494 460454 172938
rect 469794 183454 470414 218898
rect 469794 182898 469826 183454
rect 470382 182898 470414 183454
rect 461648 151174 461968 151206
rect 461648 150938 461690 151174
rect 461926 150938 461968 151174
rect 461648 150854 461968 150938
rect 461648 150618 461690 150854
rect 461926 150618 461968 150854
rect 461648 150586 461968 150618
rect 459834 136938 459866 137494
rect 460422 136938 460454 137494
rect 459834 101494 460454 136938
rect 469794 147454 470414 182898
rect 469794 146898 469826 147454
rect 470382 146898 470414 147454
rect 461648 115174 461968 115206
rect 461648 114938 461690 115174
rect 461926 114938 461968 115174
rect 461648 114854 461968 114938
rect 461648 114618 461690 114854
rect 461926 114618 461968 114854
rect 461648 114586 461968 114618
rect 459834 100938 459866 101494
rect 460422 100938 460454 101494
rect 459834 65494 460454 100938
rect 469794 111454 470414 146898
rect 469794 110898 469826 111454
rect 470382 110898 470414 111454
rect 461648 79174 461968 79206
rect 461648 78938 461690 79174
rect 461926 78938 461968 79174
rect 461648 78854 461968 78938
rect 461648 78618 461690 78854
rect 461926 78618 461968 78854
rect 461648 78586 461968 78618
rect 459834 64938 459866 65494
rect 460422 64938 460454 65494
rect 459834 29494 460454 64938
rect 469794 75454 470414 110898
rect 469794 74898 469826 75454
rect 470382 74898 470414 75454
rect 461648 43174 461968 43206
rect 461648 42938 461690 43174
rect 461926 42938 461968 43174
rect 461648 42854 461968 42938
rect 461648 42618 461690 42854
rect 461926 42618 461968 42854
rect 461648 42586 461968 42618
rect 459834 28938 459866 29494
rect 460422 28938 460454 29494
rect 459834 -7066 460454 28938
rect 469794 39454 470414 74898
rect 469794 38898 469826 39454
rect 470382 38898 470414 39454
rect 461648 7174 461968 7206
rect 461648 6938 461690 7174
rect 461926 6938 461968 7174
rect 461648 6854 461968 6938
rect 461648 6618 461690 6854
rect 461926 6618 461968 6854
rect 461648 6586 461968 6618
rect 459834 -7622 459866 -7066
rect 460422 -7622 460454 -7066
rect 459834 -7654 460454 -7622
rect 469794 3454 470414 38898
rect 469794 2898 469826 3454
rect 470382 2898 470414 3454
rect 469794 -346 470414 2898
rect 469794 -902 469826 -346
rect 470382 -902 470414 -346
rect 469794 -7654 470414 -902
rect 473514 705798 474134 711590
rect 473514 705242 473546 705798
rect 474102 705242 474134 705798
rect 473514 691174 474134 705242
rect 473514 690618 473546 691174
rect 474102 690618 474134 691174
rect 473514 655174 474134 690618
rect 473514 654618 473546 655174
rect 474102 654618 474134 655174
rect 473514 619174 474134 654618
rect 473514 618618 473546 619174
rect 474102 618618 474134 619174
rect 473514 583174 474134 618618
rect 473514 582618 473546 583174
rect 474102 582618 474134 583174
rect 473514 547174 474134 582618
rect 473514 546618 473546 547174
rect 474102 546618 474134 547174
rect 473514 511174 474134 546618
rect 473514 510618 473546 511174
rect 474102 510618 474134 511174
rect 473514 475174 474134 510618
rect 473514 474618 473546 475174
rect 474102 474618 474134 475174
rect 473514 439174 474134 474618
rect 473514 438618 473546 439174
rect 474102 438618 474134 439174
rect 473514 403174 474134 438618
rect 473514 402618 473546 403174
rect 474102 402618 474134 403174
rect 473514 367174 474134 402618
rect 473514 366618 473546 367174
rect 474102 366618 474134 367174
rect 473514 331174 474134 366618
rect 477234 706758 477854 711590
rect 477234 706202 477266 706758
rect 477822 706202 477854 706758
rect 477234 694894 477854 706202
rect 477234 694338 477266 694894
rect 477822 694338 477854 694894
rect 477234 658894 477854 694338
rect 477234 658338 477266 658894
rect 477822 658338 477854 658894
rect 477234 622894 477854 658338
rect 477234 622338 477266 622894
rect 477822 622338 477854 622894
rect 477234 586894 477854 622338
rect 477234 586338 477266 586894
rect 477822 586338 477854 586894
rect 477234 550894 477854 586338
rect 477234 550338 477266 550894
rect 477822 550338 477854 550894
rect 477234 514894 477854 550338
rect 477234 514338 477266 514894
rect 477822 514338 477854 514894
rect 477234 478894 477854 514338
rect 477234 478338 477266 478894
rect 477822 478338 477854 478894
rect 477234 442894 477854 478338
rect 477234 442338 477266 442894
rect 477822 442338 477854 442894
rect 477234 406894 477854 442338
rect 477234 406338 477266 406894
rect 477822 406338 477854 406894
rect 477234 370894 477854 406338
rect 477234 370338 477266 370894
rect 477822 370338 477854 370894
rect 477234 354900 477854 370338
rect 480954 707718 481574 711590
rect 480954 707162 480986 707718
rect 481542 707162 481574 707718
rect 480954 698614 481574 707162
rect 480954 698058 480986 698614
rect 481542 698058 481574 698614
rect 480954 662614 481574 698058
rect 480954 662058 480986 662614
rect 481542 662058 481574 662614
rect 480954 626614 481574 662058
rect 480954 626058 480986 626614
rect 481542 626058 481574 626614
rect 480954 590614 481574 626058
rect 480954 590058 480986 590614
rect 481542 590058 481574 590614
rect 480954 554614 481574 590058
rect 480954 554058 480986 554614
rect 481542 554058 481574 554614
rect 480954 518614 481574 554058
rect 480954 518058 480986 518614
rect 481542 518058 481574 518614
rect 480954 482614 481574 518058
rect 480954 482058 480986 482614
rect 481542 482058 481574 482614
rect 480954 446614 481574 482058
rect 480954 446058 480986 446614
rect 481542 446058 481574 446614
rect 480954 410614 481574 446058
rect 480954 410058 480986 410614
rect 481542 410058 481574 410614
rect 480954 374614 481574 410058
rect 480954 374058 480986 374614
rect 481542 374058 481574 374614
rect 473514 330618 473546 331174
rect 474102 330618 474134 331174
rect 473514 295174 474134 330618
rect 480954 338614 481574 374058
rect 480954 338058 480986 338614
rect 481542 338058 481574 338614
rect 477008 327454 477328 327486
rect 477008 327218 477050 327454
rect 477286 327218 477328 327454
rect 477008 327134 477328 327218
rect 477008 326898 477050 327134
rect 477286 326898 477328 327134
rect 477008 326866 477328 326898
rect 473514 294618 473546 295174
rect 474102 294618 474134 295174
rect 473514 259174 474134 294618
rect 480954 302614 481574 338058
rect 480954 302058 480986 302614
rect 481542 302058 481574 302614
rect 477008 291454 477328 291486
rect 477008 291218 477050 291454
rect 477286 291218 477328 291454
rect 477008 291134 477328 291218
rect 477008 290898 477050 291134
rect 477286 290898 477328 291134
rect 477008 290866 477328 290898
rect 473514 258618 473546 259174
rect 474102 258618 474134 259174
rect 473514 223174 474134 258618
rect 480954 266614 481574 302058
rect 480954 266058 480986 266614
rect 481542 266058 481574 266614
rect 477008 255454 477328 255486
rect 477008 255218 477050 255454
rect 477286 255218 477328 255454
rect 477008 255134 477328 255218
rect 477008 254898 477050 255134
rect 477286 254898 477328 255134
rect 477008 254866 477328 254898
rect 473514 222618 473546 223174
rect 474102 222618 474134 223174
rect 473514 187174 474134 222618
rect 480954 230614 481574 266058
rect 480954 230058 480986 230614
rect 481542 230058 481574 230614
rect 477008 219454 477328 219486
rect 477008 219218 477050 219454
rect 477286 219218 477328 219454
rect 477008 219134 477328 219218
rect 477008 218898 477050 219134
rect 477286 218898 477328 219134
rect 477008 218866 477328 218898
rect 473514 186618 473546 187174
rect 474102 186618 474134 187174
rect 473514 151174 474134 186618
rect 480954 194614 481574 230058
rect 480954 194058 480986 194614
rect 481542 194058 481574 194614
rect 477008 183454 477328 183486
rect 477008 183218 477050 183454
rect 477286 183218 477328 183454
rect 477008 183134 477328 183218
rect 477008 182898 477050 183134
rect 477286 182898 477328 183134
rect 477008 182866 477328 182898
rect 473514 150618 473546 151174
rect 474102 150618 474134 151174
rect 473514 115174 474134 150618
rect 480954 158614 481574 194058
rect 480954 158058 480986 158614
rect 481542 158058 481574 158614
rect 477008 147454 477328 147486
rect 477008 147218 477050 147454
rect 477286 147218 477328 147454
rect 477008 147134 477328 147218
rect 477008 146898 477050 147134
rect 477286 146898 477328 147134
rect 477008 146866 477328 146898
rect 473514 114618 473546 115174
rect 474102 114618 474134 115174
rect 473514 79174 474134 114618
rect 480954 122614 481574 158058
rect 480954 122058 480986 122614
rect 481542 122058 481574 122614
rect 477008 111454 477328 111486
rect 477008 111218 477050 111454
rect 477286 111218 477328 111454
rect 477008 111134 477328 111218
rect 477008 110898 477050 111134
rect 477286 110898 477328 111134
rect 477008 110866 477328 110898
rect 473514 78618 473546 79174
rect 474102 78618 474134 79174
rect 473514 43174 474134 78618
rect 480954 86614 481574 122058
rect 480954 86058 480986 86614
rect 481542 86058 481574 86614
rect 477008 75454 477328 75486
rect 477008 75218 477050 75454
rect 477286 75218 477328 75454
rect 477008 75134 477328 75218
rect 477008 74898 477050 75134
rect 477286 74898 477328 75134
rect 477008 74866 477328 74898
rect 473514 42618 473546 43174
rect 474102 42618 474134 43174
rect 473514 7174 474134 42618
rect 480954 50614 481574 86058
rect 480954 50058 480986 50614
rect 481542 50058 481574 50614
rect 477008 39454 477328 39486
rect 477008 39218 477050 39454
rect 477286 39218 477328 39454
rect 477008 39134 477328 39218
rect 477008 38898 477050 39134
rect 477286 38898 477328 39134
rect 477008 38866 477328 38898
rect 473514 6618 473546 7174
rect 474102 6618 474134 7174
rect 473514 -1306 474134 6618
rect 473514 -1862 473546 -1306
rect 474102 -1862 474134 -1306
rect 473514 -7654 474134 -1862
rect 480954 14614 481574 50058
rect 480954 14058 480986 14614
rect 481542 14058 481574 14614
rect 480954 -3226 481574 14058
rect 480954 -3782 480986 -3226
rect 481542 -3782 481574 -3226
rect 480954 -7654 481574 -3782
rect 484674 708678 485294 711590
rect 484674 708122 484706 708678
rect 485262 708122 485294 708678
rect 484674 666334 485294 708122
rect 484674 665778 484706 666334
rect 485262 665778 485294 666334
rect 484674 630334 485294 665778
rect 484674 629778 484706 630334
rect 485262 629778 485294 630334
rect 484674 594334 485294 629778
rect 484674 593778 484706 594334
rect 485262 593778 485294 594334
rect 484674 558334 485294 593778
rect 484674 557778 484706 558334
rect 485262 557778 485294 558334
rect 484674 522334 485294 557778
rect 484674 521778 484706 522334
rect 485262 521778 485294 522334
rect 484674 486334 485294 521778
rect 484674 485778 484706 486334
rect 485262 485778 485294 486334
rect 484674 450334 485294 485778
rect 484674 449778 484706 450334
rect 485262 449778 485294 450334
rect 484674 414334 485294 449778
rect 484674 413778 484706 414334
rect 485262 413778 485294 414334
rect 484674 378334 485294 413778
rect 484674 377778 484706 378334
rect 485262 377778 485294 378334
rect 484674 342334 485294 377778
rect 484674 341778 484706 342334
rect 485262 341778 485294 342334
rect 484674 306334 485294 341778
rect 484674 305778 484706 306334
rect 485262 305778 485294 306334
rect 484674 270334 485294 305778
rect 484674 269778 484706 270334
rect 485262 269778 485294 270334
rect 484674 234334 485294 269778
rect 484674 233778 484706 234334
rect 485262 233778 485294 234334
rect 484674 198334 485294 233778
rect 484674 197778 484706 198334
rect 485262 197778 485294 198334
rect 484674 162334 485294 197778
rect 484674 161778 484706 162334
rect 485262 161778 485294 162334
rect 484674 126334 485294 161778
rect 484674 125778 484706 126334
rect 485262 125778 485294 126334
rect 484674 90334 485294 125778
rect 484674 89778 484706 90334
rect 485262 89778 485294 90334
rect 484674 54334 485294 89778
rect 484674 53778 484706 54334
rect 485262 53778 485294 54334
rect 484674 18334 485294 53778
rect 484674 17778 484706 18334
rect 485262 17778 485294 18334
rect 484674 -4186 485294 17778
rect 484674 -4742 484706 -4186
rect 485262 -4742 485294 -4186
rect 484674 -7654 485294 -4742
rect 488394 709638 489014 711590
rect 488394 709082 488426 709638
rect 488982 709082 489014 709638
rect 488394 670054 489014 709082
rect 488394 669498 488426 670054
rect 488982 669498 489014 670054
rect 488394 634054 489014 669498
rect 488394 633498 488426 634054
rect 488982 633498 489014 634054
rect 488394 598054 489014 633498
rect 488394 597498 488426 598054
rect 488982 597498 489014 598054
rect 488394 562054 489014 597498
rect 488394 561498 488426 562054
rect 488982 561498 489014 562054
rect 488394 526054 489014 561498
rect 488394 525498 488426 526054
rect 488982 525498 489014 526054
rect 488394 490054 489014 525498
rect 488394 489498 488426 490054
rect 488982 489498 489014 490054
rect 488394 454054 489014 489498
rect 488394 453498 488426 454054
rect 488982 453498 489014 454054
rect 488394 418054 489014 453498
rect 488394 417498 488426 418054
rect 488982 417498 489014 418054
rect 488394 382054 489014 417498
rect 488394 381498 488426 382054
rect 488982 381498 489014 382054
rect 488394 346054 489014 381498
rect 492114 710598 492734 711590
rect 492114 710042 492146 710598
rect 492702 710042 492734 710598
rect 492114 673774 492734 710042
rect 492114 673218 492146 673774
rect 492702 673218 492734 673774
rect 492114 637774 492734 673218
rect 492114 637218 492146 637774
rect 492702 637218 492734 637774
rect 492114 601774 492734 637218
rect 492114 601218 492146 601774
rect 492702 601218 492734 601774
rect 492114 565774 492734 601218
rect 492114 565218 492146 565774
rect 492702 565218 492734 565774
rect 492114 529774 492734 565218
rect 492114 529218 492146 529774
rect 492702 529218 492734 529774
rect 492114 493774 492734 529218
rect 492114 493218 492146 493774
rect 492702 493218 492734 493774
rect 492114 457774 492734 493218
rect 492114 457218 492146 457774
rect 492702 457218 492734 457774
rect 492114 421774 492734 457218
rect 492114 421218 492146 421774
rect 492702 421218 492734 421774
rect 492114 385774 492734 421218
rect 492114 385218 492146 385774
rect 492702 385218 492734 385774
rect 492114 354900 492734 385218
rect 495834 711558 496454 711590
rect 495834 711002 495866 711558
rect 496422 711002 496454 711558
rect 495834 677494 496454 711002
rect 495834 676938 495866 677494
rect 496422 676938 496454 677494
rect 495834 641494 496454 676938
rect 495834 640938 495866 641494
rect 496422 640938 496454 641494
rect 495834 605494 496454 640938
rect 495834 604938 495866 605494
rect 496422 604938 496454 605494
rect 495834 569494 496454 604938
rect 495834 568938 495866 569494
rect 496422 568938 496454 569494
rect 495834 533494 496454 568938
rect 495834 532938 495866 533494
rect 496422 532938 496454 533494
rect 495834 497494 496454 532938
rect 495834 496938 495866 497494
rect 496422 496938 496454 497494
rect 495834 461494 496454 496938
rect 495834 460938 495866 461494
rect 496422 460938 496454 461494
rect 495834 425494 496454 460938
rect 495834 424938 495866 425494
rect 496422 424938 496454 425494
rect 495834 389494 496454 424938
rect 495834 388938 495866 389494
rect 496422 388938 496454 389494
rect 488394 345498 488426 346054
rect 488982 345498 489014 346054
rect 488394 310054 489014 345498
rect 495834 353494 496454 388938
rect 495834 352938 495866 353494
rect 496422 352938 496454 353494
rect 492368 331174 492688 331206
rect 492368 330938 492410 331174
rect 492646 330938 492688 331174
rect 492368 330854 492688 330938
rect 492368 330618 492410 330854
rect 492646 330618 492688 330854
rect 492368 330586 492688 330618
rect 488394 309498 488426 310054
rect 488982 309498 489014 310054
rect 488394 274054 489014 309498
rect 495834 317494 496454 352938
rect 495834 316938 495866 317494
rect 496422 316938 496454 317494
rect 492368 295174 492688 295206
rect 492368 294938 492410 295174
rect 492646 294938 492688 295174
rect 492368 294854 492688 294938
rect 492368 294618 492410 294854
rect 492646 294618 492688 294854
rect 492368 294586 492688 294618
rect 488394 273498 488426 274054
rect 488982 273498 489014 274054
rect 488394 238054 489014 273498
rect 495834 281494 496454 316938
rect 495834 280938 495866 281494
rect 496422 280938 496454 281494
rect 492368 259174 492688 259206
rect 492368 258938 492410 259174
rect 492646 258938 492688 259174
rect 492368 258854 492688 258938
rect 492368 258618 492410 258854
rect 492646 258618 492688 258854
rect 492368 258586 492688 258618
rect 488394 237498 488426 238054
rect 488982 237498 489014 238054
rect 488394 202054 489014 237498
rect 495834 245494 496454 280938
rect 495834 244938 495866 245494
rect 496422 244938 496454 245494
rect 492368 223174 492688 223206
rect 492368 222938 492410 223174
rect 492646 222938 492688 223174
rect 492368 222854 492688 222938
rect 492368 222618 492410 222854
rect 492646 222618 492688 222854
rect 492368 222586 492688 222618
rect 488394 201498 488426 202054
rect 488982 201498 489014 202054
rect 488394 166054 489014 201498
rect 495834 209494 496454 244938
rect 495834 208938 495866 209494
rect 496422 208938 496454 209494
rect 492368 187174 492688 187206
rect 492368 186938 492410 187174
rect 492646 186938 492688 187174
rect 492368 186854 492688 186938
rect 492368 186618 492410 186854
rect 492646 186618 492688 186854
rect 492368 186586 492688 186618
rect 488394 165498 488426 166054
rect 488982 165498 489014 166054
rect 488394 130054 489014 165498
rect 495834 173494 496454 208938
rect 495834 172938 495866 173494
rect 496422 172938 496454 173494
rect 492368 151174 492688 151206
rect 492368 150938 492410 151174
rect 492646 150938 492688 151174
rect 492368 150854 492688 150938
rect 492368 150618 492410 150854
rect 492646 150618 492688 150854
rect 492368 150586 492688 150618
rect 488394 129498 488426 130054
rect 488982 129498 489014 130054
rect 488394 94054 489014 129498
rect 495834 137494 496454 172938
rect 495834 136938 495866 137494
rect 496422 136938 496454 137494
rect 492368 115174 492688 115206
rect 492368 114938 492410 115174
rect 492646 114938 492688 115174
rect 492368 114854 492688 114938
rect 492368 114618 492410 114854
rect 492646 114618 492688 114854
rect 492368 114586 492688 114618
rect 488394 93498 488426 94054
rect 488982 93498 489014 94054
rect 488394 58054 489014 93498
rect 495834 101494 496454 136938
rect 495834 100938 495866 101494
rect 496422 100938 496454 101494
rect 492368 79174 492688 79206
rect 492368 78938 492410 79174
rect 492646 78938 492688 79174
rect 492368 78854 492688 78938
rect 492368 78618 492410 78854
rect 492646 78618 492688 78854
rect 492368 78586 492688 78618
rect 488394 57498 488426 58054
rect 488982 57498 489014 58054
rect 488394 22054 489014 57498
rect 495834 65494 496454 100938
rect 495834 64938 495866 65494
rect 496422 64938 496454 65494
rect 492368 43174 492688 43206
rect 492368 42938 492410 43174
rect 492646 42938 492688 43174
rect 492368 42854 492688 42938
rect 492368 42618 492410 42854
rect 492646 42618 492688 42854
rect 492368 42586 492688 42618
rect 488394 21498 488426 22054
rect 488982 21498 489014 22054
rect 488394 -5146 489014 21498
rect 495834 29494 496454 64938
rect 495834 28938 495866 29494
rect 496422 28938 496454 29494
rect 492368 7174 492688 7206
rect 492368 6938 492410 7174
rect 492646 6938 492688 7174
rect 492368 6854 492688 6938
rect 492368 6618 492410 6854
rect 492646 6618 492688 6854
rect 492368 6586 492688 6618
rect 488394 -5702 488426 -5146
rect 488982 -5702 489014 -5146
rect 488394 -7654 489014 -5702
rect 495834 -7066 496454 28938
rect 495834 -7622 495866 -7066
rect 496422 -7622 496454 -7066
rect 495834 -7654 496454 -7622
rect 505794 704838 506414 711590
rect 505794 704282 505826 704838
rect 506382 704282 506414 704838
rect 505794 687454 506414 704282
rect 505794 686898 505826 687454
rect 506382 686898 506414 687454
rect 505794 651454 506414 686898
rect 505794 650898 505826 651454
rect 506382 650898 506414 651454
rect 505794 615454 506414 650898
rect 505794 614898 505826 615454
rect 506382 614898 506414 615454
rect 505794 579454 506414 614898
rect 505794 578898 505826 579454
rect 506382 578898 506414 579454
rect 505794 543454 506414 578898
rect 505794 542898 505826 543454
rect 506382 542898 506414 543454
rect 505794 507454 506414 542898
rect 505794 506898 505826 507454
rect 506382 506898 506414 507454
rect 505794 471454 506414 506898
rect 505794 470898 505826 471454
rect 506382 470898 506414 471454
rect 505794 435454 506414 470898
rect 505794 434898 505826 435454
rect 506382 434898 506414 435454
rect 505794 399454 506414 434898
rect 505794 398898 505826 399454
rect 506382 398898 506414 399454
rect 505794 363454 506414 398898
rect 505794 362898 505826 363454
rect 506382 362898 506414 363454
rect 505794 327454 506414 362898
rect 509514 705798 510134 711590
rect 509514 705242 509546 705798
rect 510102 705242 510134 705798
rect 509514 691174 510134 705242
rect 509514 690618 509546 691174
rect 510102 690618 510134 691174
rect 509514 655174 510134 690618
rect 509514 654618 509546 655174
rect 510102 654618 510134 655174
rect 509514 619174 510134 654618
rect 509514 618618 509546 619174
rect 510102 618618 510134 619174
rect 509514 583174 510134 618618
rect 509514 582618 509546 583174
rect 510102 582618 510134 583174
rect 509514 547174 510134 582618
rect 509514 546618 509546 547174
rect 510102 546618 510134 547174
rect 509514 511174 510134 546618
rect 509514 510618 509546 511174
rect 510102 510618 510134 511174
rect 509514 475174 510134 510618
rect 509514 474618 509546 475174
rect 510102 474618 510134 475174
rect 509514 439174 510134 474618
rect 509514 438618 509546 439174
rect 510102 438618 510134 439174
rect 509514 403174 510134 438618
rect 509514 402618 509546 403174
rect 510102 402618 510134 403174
rect 509514 367174 510134 402618
rect 509514 366618 509546 367174
rect 510102 366618 510134 367174
rect 509514 331174 510134 366618
rect 509514 330618 509546 331174
rect 510102 330618 510134 331174
rect 505794 326898 505826 327454
rect 506382 326898 506414 327454
rect 505794 291454 506414 326898
rect 507728 327454 508048 327486
rect 507728 327218 507770 327454
rect 508006 327218 508048 327454
rect 507728 327134 508048 327218
rect 507728 326898 507770 327134
rect 508006 326898 508048 327134
rect 507728 326866 508048 326898
rect 509514 295174 510134 330618
rect 509514 294618 509546 295174
rect 510102 294618 510134 295174
rect 505794 290898 505826 291454
rect 506382 290898 506414 291454
rect 505794 255454 506414 290898
rect 507728 291454 508048 291486
rect 507728 291218 507770 291454
rect 508006 291218 508048 291454
rect 507728 291134 508048 291218
rect 507728 290898 507770 291134
rect 508006 290898 508048 291134
rect 507728 290866 508048 290898
rect 509514 259174 510134 294618
rect 509514 258618 509546 259174
rect 510102 258618 510134 259174
rect 505794 254898 505826 255454
rect 506382 254898 506414 255454
rect 505794 219454 506414 254898
rect 507728 255454 508048 255486
rect 507728 255218 507770 255454
rect 508006 255218 508048 255454
rect 507728 255134 508048 255218
rect 507728 254898 507770 255134
rect 508006 254898 508048 255134
rect 507728 254866 508048 254898
rect 509514 223174 510134 258618
rect 509514 222618 509546 223174
rect 510102 222618 510134 223174
rect 505794 218898 505826 219454
rect 506382 218898 506414 219454
rect 505794 183454 506414 218898
rect 507728 219454 508048 219486
rect 507728 219218 507770 219454
rect 508006 219218 508048 219454
rect 507728 219134 508048 219218
rect 507728 218898 507770 219134
rect 508006 218898 508048 219134
rect 507728 218866 508048 218898
rect 509514 187174 510134 222618
rect 509514 186618 509546 187174
rect 510102 186618 510134 187174
rect 505794 182898 505826 183454
rect 506382 182898 506414 183454
rect 505794 147454 506414 182898
rect 507728 183454 508048 183486
rect 507728 183218 507770 183454
rect 508006 183218 508048 183454
rect 507728 183134 508048 183218
rect 507728 182898 507770 183134
rect 508006 182898 508048 183134
rect 507728 182866 508048 182898
rect 509514 151174 510134 186618
rect 509514 150618 509546 151174
rect 510102 150618 510134 151174
rect 505794 146898 505826 147454
rect 506382 146898 506414 147454
rect 505794 111454 506414 146898
rect 507728 147454 508048 147486
rect 507728 147218 507770 147454
rect 508006 147218 508048 147454
rect 507728 147134 508048 147218
rect 507728 146898 507770 147134
rect 508006 146898 508048 147134
rect 507728 146866 508048 146898
rect 509514 115174 510134 150618
rect 509514 114618 509546 115174
rect 510102 114618 510134 115174
rect 505794 110898 505826 111454
rect 506382 110898 506414 111454
rect 505794 75454 506414 110898
rect 507728 111454 508048 111486
rect 507728 111218 507770 111454
rect 508006 111218 508048 111454
rect 507728 111134 508048 111218
rect 507728 110898 507770 111134
rect 508006 110898 508048 111134
rect 507728 110866 508048 110898
rect 509514 79174 510134 114618
rect 509514 78618 509546 79174
rect 510102 78618 510134 79174
rect 505794 74898 505826 75454
rect 506382 74898 506414 75454
rect 505794 39454 506414 74898
rect 507728 75454 508048 75486
rect 507728 75218 507770 75454
rect 508006 75218 508048 75454
rect 507728 75134 508048 75218
rect 507728 74898 507770 75134
rect 508006 74898 508048 75134
rect 507728 74866 508048 74898
rect 509514 43174 510134 78618
rect 509514 42618 509546 43174
rect 510102 42618 510134 43174
rect 505794 38898 505826 39454
rect 506382 38898 506414 39454
rect 505794 3454 506414 38898
rect 507728 39454 508048 39486
rect 507728 39218 507770 39454
rect 508006 39218 508048 39454
rect 507728 39134 508048 39218
rect 507728 38898 507770 39134
rect 508006 38898 508048 39134
rect 507728 38866 508048 38898
rect 505794 2898 505826 3454
rect 506382 2898 506414 3454
rect 505794 -346 506414 2898
rect 505794 -902 505826 -346
rect 506382 -902 506414 -346
rect 505794 -7654 506414 -902
rect 509514 7174 510134 42618
rect 509514 6618 509546 7174
rect 510102 6618 510134 7174
rect 509514 -1306 510134 6618
rect 509514 -1862 509546 -1306
rect 510102 -1862 510134 -1306
rect 509514 -7654 510134 -1862
rect 513234 706758 513854 711590
rect 513234 706202 513266 706758
rect 513822 706202 513854 706758
rect 513234 694894 513854 706202
rect 513234 694338 513266 694894
rect 513822 694338 513854 694894
rect 513234 658894 513854 694338
rect 513234 658338 513266 658894
rect 513822 658338 513854 658894
rect 513234 622894 513854 658338
rect 513234 622338 513266 622894
rect 513822 622338 513854 622894
rect 513234 586894 513854 622338
rect 513234 586338 513266 586894
rect 513822 586338 513854 586894
rect 513234 550894 513854 586338
rect 513234 550338 513266 550894
rect 513822 550338 513854 550894
rect 513234 514894 513854 550338
rect 513234 514338 513266 514894
rect 513822 514338 513854 514894
rect 513234 478894 513854 514338
rect 513234 478338 513266 478894
rect 513822 478338 513854 478894
rect 513234 442894 513854 478338
rect 513234 442338 513266 442894
rect 513822 442338 513854 442894
rect 513234 406894 513854 442338
rect 513234 406338 513266 406894
rect 513822 406338 513854 406894
rect 513234 370894 513854 406338
rect 513234 370338 513266 370894
rect 513822 370338 513854 370894
rect 513234 334894 513854 370338
rect 513234 334338 513266 334894
rect 513822 334338 513854 334894
rect 513234 298894 513854 334338
rect 513234 298338 513266 298894
rect 513822 298338 513854 298894
rect 513234 262894 513854 298338
rect 513234 262338 513266 262894
rect 513822 262338 513854 262894
rect 513234 226894 513854 262338
rect 513234 226338 513266 226894
rect 513822 226338 513854 226894
rect 513234 190894 513854 226338
rect 513234 190338 513266 190894
rect 513822 190338 513854 190894
rect 513234 154894 513854 190338
rect 513234 154338 513266 154894
rect 513822 154338 513854 154894
rect 513234 118894 513854 154338
rect 513234 118338 513266 118894
rect 513822 118338 513854 118894
rect 513234 82894 513854 118338
rect 513234 82338 513266 82894
rect 513822 82338 513854 82894
rect 513234 46894 513854 82338
rect 513234 46338 513266 46894
rect 513822 46338 513854 46894
rect 513234 10894 513854 46338
rect 513234 10338 513266 10894
rect 513822 10338 513854 10894
rect 513234 -2266 513854 10338
rect 513234 -2822 513266 -2266
rect 513822 -2822 513854 -2266
rect 513234 -7654 513854 -2822
rect 516954 707718 517574 711590
rect 516954 707162 516986 707718
rect 517542 707162 517574 707718
rect 516954 698614 517574 707162
rect 516954 698058 516986 698614
rect 517542 698058 517574 698614
rect 516954 662614 517574 698058
rect 516954 662058 516986 662614
rect 517542 662058 517574 662614
rect 516954 626614 517574 662058
rect 516954 626058 516986 626614
rect 517542 626058 517574 626614
rect 516954 590614 517574 626058
rect 516954 590058 516986 590614
rect 517542 590058 517574 590614
rect 516954 554614 517574 590058
rect 516954 554058 516986 554614
rect 517542 554058 517574 554614
rect 516954 518614 517574 554058
rect 516954 518058 516986 518614
rect 517542 518058 517574 518614
rect 516954 482614 517574 518058
rect 516954 482058 516986 482614
rect 517542 482058 517574 482614
rect 516954 446614 517574 482058
rect 516954 446058 516986 446614
rect 517542 446058 517574 446614
rect 516954 410614 517574 446058
rect 516954 410058 516986 410614
rect 517542 410058 517574 410614
rect 516954 374614 517574 410058
rect 516954 374058 516986 374614
rect 517542 374058 517574 374614
rect 516954 338614 517574 374058
rect 516954 338058 516986 338614
rect 517542 338058 517574 338614
rect 516954 302614 517574 338058
rect 516954 302058 516986 302614
rect 517542 302058 517574 302614
rect 516954 266614 517574 302058
rect 516954 266058 516986 266614
rect 517542 266058 517574 266614
rect 516954 230614 517574 266058
rect 516954 230058 516986 230614
rect 517542 230058 517574 230614
rect 516954 194614 517574 230058
rect 516954 194058 516986 194614
rect 517542 194058 517574 194614
rect 516954 158614 517574 194058
rect 516954 158058 516986 158614
rect 517542 158058 517574 158614
rect 516954 122614 517574 158058
rect 516954 122058 516986 122614
rect 517542 122058 517574 122614
rect 516954 86614 517574 122058
rect 516954 86058 516986 86614
rect 517542 86058 517574 86614
rect 516954 50614 517574 86058
rect 516954 50058 516986 50614
rect 517542 50058 517574 50614
rect 516954 14614 517574 50058
rect 516954 14058 516986 14614
rect 517542 14058 517574 14614
rect 516954 -3226 517574 14058
rect 516954 -3782 516986 -3226
rect 517542 -3782 517574 -3226
rect 516954 -7654 517574 -3782
rect 520674 708678 521294 711590
rect 520674 708122 520706 708678
rect 521262 708122 521294 708678
rect 520674 666334 521294 708122
rect 520674 665778 520706 666334
rect 521262 665778 521294 666334
rect 520674 630334 521294 665778
rect 520674 629778 520706 630334
rect 521262 629778 521294 630334
rect 520674 594334 521294 629778
rect 520674 593778 520706 594334
rect 521262 593778 521294 594334
rect 520674 558334 521294 593778
rect 520674 557778 520706 558334
rect 521262 557778 521294 558334
rect 520674 522334 521294 557778
rect 520674 521778 520706 522334
rect 521262 521778 521294 522334
rect 520674 486334 521294 521778
rect 520674 485778 520706 486334
rect 521262 485778 521294 486334
rect 520674 450334 521294 485778
rect 520674 449778 520706 450334
rect 521262 449778 521294 450334
rect 520674 414334 521294 449778
rect 520674 413778 520706 414334
rect 521262 413778 521294 414334
rect 520674 378334 521294 413778
rect 520674 377778 520706 378334
rect 521262 377778 521294 378334
rect 520674 342334 521294 377778
rect 520674 341778 520706 342334
rect 521262 341778 521294 342334
rect 520674 306334 521294 341778
rect 524394 709638 525014 711590
rect 524394 709082 524426 709638
rect 524982 709082 525014 709638
rect 524394 670054 525014 709082
rect 524394 669498 524426 670054
rect 524982 669498 525014 670054
rect 524394 634054 525014 669498
rect 524394 633498 524426 634054
rect 524982 633498 525014 634054
rect 524394 598054 525014 633498
rect 524394 597498 524426 598054
rect 524982 597498 525014 598054
rect 524394 562054 525014 597498
rect 524394 561498 524426 562054
rect 524982 561498 525014 562054
rect 524394 526054 525014 561498
rect 524394 525498 524426 526054
rect 524982 525498 525014 526054
rect 524394 490054 525014 525498
rect 524394 489498 524426 490054
rect 524982 489498 525014 490054
rect 524394 454054 525014 489498
rect 524394 453498 524426 454054
rect 524982 453498 525014 454054
rect 524394 418054 525014 453498
rect 524394 417498 524426 418054
rect 524982 417498 525014 418054
rect 524394 382054 525014 417498
rect 524394 381498 524426 382054
rect 524982 381498 525014 382054
rect 524394 346054 525014 381498
rect 524394 345498 524426 346054
rect 524982 345498 525014 346054
rect 523088 331174 523408 331206
rect 523088 330938 523130 331174
rect 523366 330938 523408 331174
rect 523088 330854 523408 330938
rect 523088 330618 523130 330854
rect 523366 330618 523408 330854
rect 523088 330586 523408 330618
rect 520674 305778 520706 306334
rect 521262 305778 521294 306334
rect 520674 270334 521294 305778
rect 524394 310054 525014 345498
rect 524394 309498 524426 310054
rect 524982 309498 525014 310054
rect 523088 295174 523408 295206
rect 523088 294938 523130 295174
rect 523366 294938 523408 295174
rect 523088 294854 523408 294938
rect 523088 294618 523130 294854
rect 523366 294618 523408 294854
rect 523088 294586 523408 294618
rect 520674 269778 520706 270334
rect 521262 269778 521294 270334
rect 520674 234334 521294 269778
rect 524394 274054 525014 309498
rect 524394 273498 524426 274054
rect 524982 273498 525014 274054
rect 523088 259174 523408 259206
rect 523088 258938 523130 259174
rect 523366 258938 523408 259174
rect 523088 258854 523408 258938
rect 523088 258618 523130 258854
rect 523366 258618 523408 258854
rect 523088 258586 523408 258618
rect 520674 233778 520706 234334
rect 521262 233778 521294 234334
rect 520674 198334 521294 233778
rect 524394 238054 525014 273498
rect 524394 237498 524426 238054
rect 524982 237498 525014 238054
rect 523088 223174 523408 223206
rect 523088 222938 523130 223174
rect 523366 222938 523408 223174
rect 523088 222854 523408 222938
rect 523088 222618 523130 222854
rect 523366 222618 523408 222854
rect 523088 222586 523408 222618
rect 520674 197778 520706 198334
rect 521262 197778 521294 198334
rect 520674 162334 521294 197778
rect 524394 202054 525014 237498
rect 524394 201498 524426 202054
rect 524982 201498 525014 202054
rect 523088 187174 523408 187206
rect 523088 186938 523130 187174
rect 523366 186938 523408 187174
rect 523088 186854 523408 186938
rect 523088 186618 523130 186854
rect 523366 186618 523408 186854
rect 523088 186586 523408 186618
rect 520674 161778 520706 162334
rect 521262 161778 521294 162334
rect 520674 126334 521294 161778
rect 524394 166054 525014 201498
rect 524394 165498 524426 166054
rect 524982 165498 525014 166054
rect 523088 151174 523408 151206
rect 523088 150938 523130 151174
rect 523366 150938 523408 151174
rect 523088 150854 523408 150938
rect 523088 150618 523130 150854
rect 523366 150618 523408 150854
rect 523088 150586 523408 150618
rect 520674 125778 520706 126334
rect 521262 125778 521294 126334
rect 520674 90334 521294 125778
rect 524394 130054 525014 165498
rect 524394 129498 524426 130054
rect 524982 129498 525014 130054
rect 523088 115174 523408 115206
rect 523088 114938 523130 115174
rect 523366 114938 523408 115174
rect 523088 114854 523408 114938
rect 523088 114618 523130 114854
rect 523366 114618 523408 114854
rect 523088 114586 523408 114618
rect 520674 89778 520706 90334
rect 521262 89778 521294 90334
rect 520674 54334 521294 89778
rect 524394 94054 525014 129498
rect 524394 93498 524426 94054
rect 524982 93498 525014 94054
rect 523088 79174 523408 79206
rect 523088 78938 523130 79174
rect 523366 78938 523408 79174
rect 523088 78854 523408 78938
rect 523088 78618 523130 78854
rect 523366 78618 523408 78854
rect 523088 78586 523408 78618
rect 520674 53778 520706 54334
rect 521262 53778 521294 54334
rect 520674 18334 521294 53778
rect 524394 58054 525014 93498
rect 524394 57498 524426 58054
rect 524982 57498 525014 58054
rect 523088 43174 523408 43206
rect 523088 42938 523130 43174
rect 523366 42938 523408 43174
rect 523088 42854 523408 42938
rect 523088 42618 523130 42854
rect 523366 42618 523408 42854
rect 523088 42586 523408 42618
rect 520674 17778 520706 18334
rect 521262 17778 521294 18334
rect 520674 -4186 521294 17778
rect 524394 22054 525014 57498
rect 524394 21498 524426 22054
rect 524982 21498 525014 22054
rect 523088 7174 523408 7206
rect 523088 6938 523130 7174
rect 523366 6938 523408 7174
rect 523088 6854 523408 6938
rect 523088 6618 523130 6854
rect 523366 6618 523408 6854
rect 523088 6586 523408 6618
rect 520674 -4742 520706 -4186
rect 521262 -4742 521294 -4186
rect 520674 -7654 521294 -4742
rect 524394 -5146 525014 21498
rect 524394 -5702 524426 -5146
rect 524982 -5702 525014 -5146
rect 524394 -7654 525014 -5702
rect 528114 710598 528734 711590
rect 528114 710042 528146 710598
rect 528702 710042 528734 710598
rect 528114 673774 528734 710042
rect 528114 673218 528146 673774
rect 528702 673218 528734 673774
rect 528114 637774 528734 673218
rect 528114 637218 528146 637774
rect 528702 637218 528734 637774
rect 528114 601774 528734 637218
rect 528114 601218 528146 601774
rect 528702 601218 528734 601774
rect 528114 565774 528734 601218
rect 528114 565218 528146 565774
rect 528702 565218 528734 565774
rect 528114 529774 528734 565218
rect 528114 529218 528146 529774
rect 528702 529218 528734 529774
rect 528114 493774 528734 529218
rect 528114 493218 528146 493774
rect 528702 493218 528734 493774
rect 528114 457774 528734 493218
rect 528114 457218 528146 457774
rect 528702 457218 528734 457774
rect 528114 421774 528734 457218
rect 528114 421218 528146 421774
rect 528702 421218 528734 421774
rect 528114 385774 528734 421218
rect 528114 385218 528146 385774
rect 528702 385218 528734 385774
rect 528114 349774 528734 385218
rect 528114 349218 528146 349774
rect 528702 349218 528734 349774
rect 528114 313774 528734 349218
rect 528114 313218 528146 313774
rect 528702 313218 528734 313774
rect 528114 277774 528734 313218
rect 528114 277218 528146 277774
rect 528702 277218 528734 277774
rect 528114 241774 528734 277218
rect 528114 241218 528146 241774
rect 528702 241218 528734 241774
rect 528114 205774 528734 241218
rect 528114 205218 528146 205774
rect 528702 205218 528734 205774
rect 528114 169774 528734 205218
rect 528114 169218 528146 169774
rect 528702 169218 528734 169774
rect 528114 133774 528734 169218
rect 528114 133218 528146 133774
rect 528702 133218 528734 133774
rect 528114 97774 528734 133218
rect 528114 97218 528146 97774
rect 528702 97218 528734 97774
rect 528114 61774 528734 97218
rect 528114 61218 528146 61774
rect 528702 61218 528734 61774
rect 528114 25774 528734 61218
rect 528114 25218 528146 25774
rect 528702 25218 528734 25774
rect 528114 -6106 528734 25218
rect 528114 -6662 528146 -6106
rect 528702 -6662 528734 -6106
rect 528114 -7654 528734 -6662
rect 531834 711558 532454 711590
rect 531834 711002 531866 711558
rect 532422 711002 532454 711558
rect 531834 677494 532454 711002
rect 531834 676938 531866 677494
rect 532422 676938 532454 677494
rect 531834 641494 532454 676938
rect 531834 640938 531866 641494
rect 532422 640938 532454 641494
rect 531834 605494 532454 640938
rect 531834 604938 531866 605494
rect 532422 604938 532454 605494
rect 531834 569494 532454 604938
rect 531834 568938 531866 569494
rect 532422 568938 532454 569494
rect 531834 533494 532454 568938
rect 531834 532938 531866 533494
rect 532422 532938 532454 533494
rect 531834 497494 532454 532938
rect 531834 496938 531866 497494
rect 532422 496938 532454 497494
rect 531834 461494 532454 496938
rect 531834 460938 531866 461494
rect 532422 460938 532454 461494
rect 531834 425494 532454 460938
rect 531834 424938 531866 425494
rect 532422 424938 532454 425494
rect 531834 389494 532454 424938
rect 531834 388938 531866 389494
rect 532422 388938 532454 389494
rect 531834 353494 532454 388938
rect 531834 352938 531866 353494
rect 532422 352938 532454 353494
rect 531834 317494 532454 352938
rect 541794 704838 542414 711590
rect 541794 704282 541826 704838
rect 542382 704282 542414 704838
rect 541794 687454 542414 704282
rect 541794 686898 541826 687454
rect 542382 686898 542414 687454
rect 541794 651454 542414 686898
rect 541794 650898 541826 651454
rect 542382 650898 542414 651454
rect 541794 615454 542414 650898
rect 541794 614898 541826 615454
rect 542382 614898 542414 615454
rect 541794 579454 542414 614898
rect 541794 578898 541826 579454
rect 542382 578898 542414 579454
rect 541794 543454 542414 578898
rect 541794 542898 541826 543454
rect 542382 542898 542414 543454
rect 541794 507454 542414 542898
rect 541794 506898 541826 507454
rect 542382 506898 542414 507454
rect 541794 471454 542414 506898
rect 541794 470898 541826 471454
rect 542382 470898 542414 471454
rect 541794 435454 542414 470898
rect 541794 434898 541826 435454
rect 542382 434898 542414 435454
rect 541794 399454 542414 434898
rect 541794 398898 541826 399454
rect 542382 398898 542414 399454
rect 541794 363454 542414 398898
rect 541794 362898 541826 363454
rect 542382 362898 542414 363454
rect 538448 327454 538768 327486
rect 538448 327218 538490 327454
rect 538726 327218 538768 327454
rect 538448 327134 538768 327218
rect 538448 326898 538490 327134
rect 538726 326898 538768 327134
rect 538448 326866 538768 326898
rect 541794 327454 542414 362898
rect 541794 326898 541826 327454
rect 542382 326898 542414 327454
rect 531834 316938 531866 317494
rect 532422 316938 532454 317494
rect 531834 281494 532454 316938
rect 538448 291454 538768 291486
rect 538448 291218 538490 291454
rect 538726 291218 538768 291454
rect 538448 291134 538768 291218
rect 538448 290898 538490 291134
rect 538726 290898 538768 291134
rect 538448 290866 538768 290898
rect 541794 291454 542414 326898
rect 541794 290898 541826 291454
rect 542382 290898 542414 291454
rect 531834 280938 531866 281494
rect 532422 280938 532454 281494
rect 531834 245494 532454 280938
rect 538448 255454 538768 255486
rect 538448 255218 538490 255454
rect 538726 255218 538768 255454
rect 538448 255134 538768 255218
rect 538448 254898 538490 255134
rect 538726 254898 538768 255134
rect 538448 254866 538768 254898
rect 541794 255454 542414 290898
rect 541794 254898 541826 255454
rect 542382 254898 542414 255454
rect 531834 244938 531866 245494
rect 532422 244938 532454 245494
rect 531834 209494 532454 244938
rect 538448 219454 538768 219486
rect 538448 219218 538490 219454
rect 538726 219218 538768 219454
rect 538448 219134 538768 219218
rect 538448 218898 538490 219134
rect 538726 218898 538768 219134
rect 538448 218866 538768 218898
rect 541794 219454 542414 254898
rect 541794 218898 541826 219454
rect 542382 218898 542414 219454
rect 531834 208938 531866 209494
rect 532422 208938 532454 209494
rect 531834 173494 532454 208938
rect 538448 183454 538768 183486
rect 538448 183218 538490 183454
rect 538726 183218 538768 183454
rect 538448 183134 538768 183218
rect 538448 182898 538490 183134
rect 538726 182898 538768 183134
rect 538448 182866 538768 182898
rect 541794 183454 542414 218898
rect 541794 182898 541826 183454
rect 542382 182898 542414 183454
rect 531834 172938 531866 173494
rect 532422 172938 532454 173494
rect 531834 137494 532454 172938
rect 538448 147454 538768 147486
rect 538448 147218 538490 147454
rect 538726 147218 538768 147454
rect 538448 147134 538768 147218
rect 538448 146898 538490 147134
rect 538726 146898 538768 147134
rect 538448 146866 538768 146898
rect 541794 147454 542414 182898
rect 541794 146898 541826 147454
rect 542382 146898 542414 147454
rect 531834 136938 531866 137494
rect 532422 136938 532454 137494
rect 531834 101494 532454 136938
rect 538448 111454 538768 111486
rect 538448 111218 538490 111454
rect 538726 111218 538768 111454
rect 538448 111134 538768 111218
rect 538448 110898 538490 111134
rect 538726 110898 538768 111134
rect 538448 110866 538768 110898
rect 541794 111454 542414 146898
rect 541794 110898 541826 111454
rect 542382 110898 542414 111454
rect 531834 100938 531866 101494
rect 532422 100938 532454 101494
rect 531834 65494 532454 100938
rect 538448 75454 538768 75486
rect 538448 75218 538490 75454
rect 538726 75218 538768 75454
rect 538448 75134 538768 75218
rect 538448 74898 538490 75134
rect 538726 74898 538768 75134
rect 538448 74866 538768 74898
rect 541794 75454 542414 110898
rect 541794 74898 541826 75454
rect 542382 74898 542414 75454
rect 531834 64938 531866 65494
rect 532422 64938 532454 65494
rect 531834 29494 532454 64938
rect 538448 39454 538768 39486
rect 538448 39218 538490 39454
rect 538726 39218 538768 39454
rect 538448 39134 538768 39218
rect 538448 38898 538490 39134
rect 538726 38898 538768 39134
rect 538448 38866 538768 38898
rect 541794 39454 542414 74898
rect 541794 38898 541826 39454
rect 542382 38898 542414 39454
rect 531834 28938 531866 29494
rect 532422 28938 532454 29494
rect 531834 -7066 532454 28938
rect 531834 -7622 531866 -7066
rect 532422 -7622 532454 -7066
rect 531834 -7654 532454 -7622
rect 541794 3454 542414 38898
rect 541794 2898 541826 3454
rect 542382 2898 542414 3454
rect 541794 -346 542414 2898
rect 541794 -902 541826 -346
rect 542382 -902 542414 -346
rect 541794 -7654 542414 -902
rect 545514 705798 546134 711590
rect 545514 705242 545546 705798
rect 546102 705242 546134 705798
rect 545514 691174 546134 705242
rect 545514 690618 545546 691174
rect 546102 690618 546134 691174
rect 545514 655174 546134 690618
rect 545514 654618 545546 655174
rect 546102 654618 546134 655174
rect 545514 619174 546134 654618
rect 545514 618618 545546 619174
rect 546102 618618 546134 619174
rect 545514 583174 546134 618618
rect 545514 582618 545546 583174
rect 546102 582618 546134 583174
rect 545514 547174 546134 582618
rect 545514 546618 545546 547174
rect 546102 546618 546134 547174
rect 545514 511174 546134 546618
rect 545514 510618 545546 511174
rect 546102 510618 546134 511174
rect 545514 475174 546134 510618
rect 545514 474618 545546 475174
rect 546102 474618 546134 475174
rect 545514 439174 546134 474618
rect 545514 438618 545546 439174
rect 546102 438618 546134 439174
rect 545514 403174 546134 438618
rect 545514 402618 545546 403174
rect 546102 402618 546134 403174
rect 545514 367174 546134 402618
rect 545514 366618 545546 367174
rect 546102 366618 546134 367174
rect 545514 331174 546134 366618
rect 545514 330618 545546 331174
rect 546102 330618 546134 331174
rect 545514 295174 546134 330618
rect 545514 294618 545546 295174
rect 546102 294618 546134 295174
rect 545514 259174 546134 294618
rect 545514 258618 545546 259174
rect 546102 258618 546134 259174
rect 545514 223174 546134 258618
rect 545514 222618 545546 223174
rect 546102 222618 546134 223174
rect 545514 187174 546134 222618
rect 545514 186618 545546 187174
rect 546102 186618 546134 187174
rect 545514 151174 546134 186618
rect 545514 150618 545546 151174
rect 546102 150618 546134 151174
rect 545514 115174 546134 150618
rect 545514 114618 545546 115174
rect 546102 114618 546134 115174
rect 545514 79174 546134 114618
rect 545514 78618 545546 79174
rect 546102 78618 546134 79174
rect 545514 43174 546134 78618
rect 545514 42618 545546 43174
rect 546102 42618 546134 43174
rect 545514 7174 546134 42618
rect 545514 6618 545546 7174
rect 546102 6618 546134 7174
rect 545514 -1306 546134 6618
rect 545514 -1862 545546 -1306
rect 546102 -1862 546134 -1306
rect 545514 -7654 546134 -1862
rect 549234 706758 549854 711590
rect 549234 706202 549266 706758
rect 549822 706202 549854 706758
rect 549234 694894 549854 706202
rect 549234 694338 549266 694894
rect 549822 694338 549854 694894
rect 549234 658894 549854 694338
rect 549234 658338 549266 658894
rect 549822 658338 549854 658894
rect 549234 622894 549854 658338
rect 549234 622338 549266 622894
rect 549822 622338 549854 622894
rect 549234 586894 549854 622338
rect 549234 586338 549266 586894
rect 549822 586338 549854 586894
rect 549234 550894 549854 586338
rect 549234 550338 549266 550894
rect 549822 550338 549854 550894
rect 549234 514894 549854 550338
rect 549234 514338 549266 514894
rect 549822 514338 549854 514894
rect 549234 478894 549854 514338
rect 549234 478338 549266 478894
rect 549822 478338 549854 478894
rect 549234 442894 549854 478338
rect 549234 442338 549266 442894
rect 549822 442338 549854 442894
rect 549234 406894 549854 442338
rect 549234 406338 549266 406894
rect 549822 406338 549854 406894
rect 549234 370894 549854 406338
rect 549234 370338 549266 370894
rect 549822 370338 549854 370894
rect 549234 334894 549854 370338
rect 549234 334338 549266 334894
rect 549822 334338 549854 334894
rect 549234 298894 549854 334338
rect 549234 298338 549266 298894
rect 549822 298338 549854 298894
rect 549234 262894 549854 298338
rect 549234 262338 549266 262894
rect 549822 262338 549854 262894
rect 549234 226894 549854 262338
rect 549234 226338 549266 226894
rect 549822 226338 549854 226894
rect 549234 190894 549854 226338
rect 549234 190338 549266 190894
rect 549822 190338 549854 190894
rect 549234 154894 549854 190338
rect 549234 154338 549266 154894
rect 549822 154338 549854 154894
rect 549234 118894 549854 154338
rect 549234 118338 549266 118894
rect 549822 118338 549854 118894
rect 549234 82894 549854 118338
rect 549234 82338 549266 82894
rect 549822 82338 549854 82894
rect 549234 46894 549854 82338
rect 549234 46338 549266 46894
rect 549822 46338 549854 46894
rect 549234 10894 549854 46338
rect 549234 10338 549266 10894
rect 549822 10338 549854 10894
rect 549234 -2266 549854 10338
rect 549234 -2822 549266 -2266
rect 549822 -2822 549854 -2266
rect 549234 -7654 549854 -2822
rect 552954 707718 553574 711590
rect 552954 707162 552986 707718
rect 553542 707162 553574 707718
rect 552954 698614 553574 707162
rect 552954 698058 552986 698614
rect 553542 698058 553574 698614
rect 552954 662614 553574 698058
rect 552954 662058 552986 662614
rect 553542 662058 553574 662614
rect 552954 626614 553574 662058
rect 552954 626058 552986 626614
rect 553542 626058 553574 626614
rect 552954 590614 553574 626058
rect 552954 590058 552986 590614
rect 553542 590058 553574 590614
rect 552954 554614 553574 590058
rect 552954 554058 552986 554614
rect 553542 554058 553574 554614
rect 552954 518614 553574 554058
rect 552954 518058 552986 518614
rect 553542 518058 553574 518614
rect 552954 482614 553574 518058
rect 552954 482058 552986 482614
rect 553542 482058 553574 482614
rect 552954 446614 553574 482058
rect 552954 446058 552986 446614
rect 553542 446058 553574 446614
rect 552954 410614 553574 446058
rect 552954 410058 552986 410614
rect 553542 410058 553574 410614
rect 552954 374614 553574 410058
rect 552954 374058 552986 374614
rect 553542 374058 553574 374614
rect 552954 338614 553574 374058
rect 552954 338058 552986 338614
rect 553542 338058 553574 338614
rect 552954 302614 553574 338058
rect 556674 708678 557294 711590
rect 556674 708122 556706 708678
rect 557262 708122 557294 708678
rect 556674 666334 557294 708122
rect 556674 665778 556706 666334
rect 557262 665778 557294 666334
rect 556674 630334 557294 665778
rect 556674 629778 556706 630334
rect 557262 629778 557294 630334
rect 556674 594334 557294 629778
rect 556674 593778 556706 594334
rect 557262 593778 557294 594334
rect 556674 558334 557294 593778
rect 556674 557778 556706 558334
rect 557262 557778 557294 558334
rect 556674 522334 557294 557778
rect 556674 521778 556706 522334
rect 557262 521778 557294 522334
rect 556674 486334 557294 521778
rect 556674 485778 556706 486334
rect 557262 485778 557294 486334
rect 556674 450334 557294 485778
rect 556674 449778 556706 450334
rect 557262 449778 557294 450334
rect 556674 414334 557294 449778
rect 556674 413778 556706 414334
rect 557262 413778 557294 414334
rect 556674 378334 557294 413778
rect 556674 377778 556706 378334
rect 557262 377778 557294 378334
rect 556674 342334 557294 377778
rect 556674 341778 556706 342334
rect 557262 341778 557294 342334
rect 553808 331174 554128 331206
rect 553808 330938 553850 331174
rect 554086 330938 554128 331174
rect 553808 330854 554128 330938
rect 553808 330618 553850 330854
rect 554086 330618 554128 330854
rect 553808 330586 554128 330618
rect 552954 302058 552986 302614
rect 553542 302058 553574 302614
rect 552954 266614 553574 302058
rect 556674 306334 557294 341778
rect 556674 305778 556706 306334
rect 557262 305778 557294 306334
rect 553808 295174 554128 295206
rect 553808 294938 553850 295174
rect 554086 294938 554128 295174
rect 553808 294854 554128 294938
rect 553808 294618 553850 294854
rect 554086 294618 554128 294854
rect 553808 294586 554128 294618
rect 552954 266058 552986 266614
rect 553542 266058 553574 266614
rect 552954 230614 553574 266058
rect 556674 270334 557294 305778
rect 556674 269778 556706 270334
rect 557262 269778 557294 270334
rect 553808 259174 554128 259206
rect 553808 258938 553850 259174
rect 554086 258938 554128 259174
rect 553808 258854 554128 258938
rect 553808 258618 553850 258854
rect 554086 258618 554128 258854
rect 553808 258586 554128 258618
rect 552954 230058 552986 230614
rect 553542 230058 553574 230614
rect 552954 194614 553574 230058
rect 556674 234334 557294 269778
rect 556674 233778 556706 234334
rect 557262 233778 557294 234334
rect 553808 223174 554128 223206
rect 553808 222938 553850 223174
rect 554086 222938 554128 223174
rect 553808 222854 554128 222938
rect 553808 222618 553850 222854
rect 554086 222618 554128 222854
rect 553808 222586 554128 222618
rect 552954 194058 552986 194614
rect 553542 194058 553574 194614
rect 552954 158614 553574 194058
rect 556674 198334 557294 233778
rect 556674 197778 556706 198334
rect 557262 197778 557294 198334
rect 553808 187174 554128 187206
rect 553808 186938 553850 187174
rect 554086 186938 554128 187174
rect 553808 186854 554128 186938
rect 553808 186618 553850 186854
rect 554086 186618 554128 186854
rect 553808 186586 554128 186618
rect 552954 158058 552986 158614
rect 553542 158058 553574 158614
rect 552954 122614 553574 158058
rect 556674 162334 557294 197778
rect 556674 161778 556706 162334
rect 557262 161778 557294 162334
rect 553808 151174 554128 151206
rect 553808 150938 553850 151174
rect 554086 150938 554128 151174
rect 553808 150854 554128 150938
rect 553808 150618 553850 150854
rect 554086 150618 554128 150854
rect 553808 150586 554128 150618
rect 552954 122058 552986 122614
rect 553542 122058 553574 122614
rect 552954 86614 553574 122058
rect 556674 126334 557294 161778
rect 556674 125778 556706 126334
rect 557262 125778 557294 126334
rect 553808 115174 554128 115206
rect 553808 114938 553850 115174
rect 554086 114938 554128 115174
rect 553808 114854 554128 114938
rect 553808 114618 553850 114854
rect 554086 114618 554128 114854
rect 553808 114586 554128 114618
rect 552954 86058 552986 86614
rect 553542 86058 553574 86614
rect 552954 50614 553574 86058
rect 556674 90334 557294 125778
rect 556674 89778 556706 90334
rect 557262 89778 557294 90334
rect 553808 79174 554128 79206
rect 553808 78938 553850 79174
rect 554086 78938 554128 79174
rect 553808 78854 554128 78938
rect 553808 78618 553850 78854
rect 554086 78618 554128 78854
rect 553808 78586 554128 78618
rect 552954 50058 552986 50614
rect 553542 50058 553574 50614
rect 552954 14614 553574 50058
rect 556674 54334 557294 89778
rect 556674 53778 556706 54334
rect 557262 53778 557294 54334
rect 553808 43174 554128 43206
rect 553808 42938 553850 43174
rect 554086 42938 554128 43174
rect 553808 42854 554128 42938
rect 553808 42618 553850 42854
rect 554086 42618 554128 42854
rect 553808 42586 554128 42618
rect 552954 14058 552986 14614
rect 553542 14058 553574 14614
rect 552954 -3226 553574 14058
rect 556674 18334 557294 53778
rect 556674 17778 556706 18334
rect 557262 17778 557294 18334
rect 553808 7174 554128 7206
rect 553808 6938 553850 7174
rect 554086 6938 554128 7174
rect 553808 6854 554128 6938
rect 553808 6618 553850 6854
rect 554086 6618 554128 6854
rect 553808 6586 554128 6618
rect 552954 -3782 552986 -3226
rect 553542 -3782 553574 -3226
rect 552954 -7654 553574 -3782
rect 556674 -4186 557294 17778
rect 556674 -4742 556706 -4186
rect 557262 -4742 557294 -4186
rect 556674 -7654 557294 -4742
rect 560394 709638 561014 711590
rect 560394 709082 560426 709638
rect 560982 709082 561014 709638
rect 560394 670054 561014 709082
rect 560394 669498 560426 670054
rect 560982 669498 561014 670054
rect 560394 634054 561014 669498
rect 560394 633498 560426 634054
rect 560982 633498 561014 634054
rect 560394 598054 561014 633498
rect 560394 597498 560426 598054
rect 560982 597498 561014 598054
rect 560394 562054 561014 597498
rect 560394 561498 560426 562054
rect 560982 561498 561014 562054
rect 560394 526054 561014 561498
rect 560394 525498 560426 526054
rect 560982 525498 561014 526054
rect 560394 490054 561014 525498
rect 560394 489498 560426 490054
rect 560982 489498 561014 490054
rect 560394 454054 561014 489498
rect 560394 453498 560426 454054
rect 560982 453498 561014 454054
rect 560394 418054 561014 453498
rect 560394 417498 560426 418054
rect 560982 417498 561014 418054
rect 560394 382054 561014 417498
rect 560394 381498 560426 382054
rect 560982 381498 561014 382054
rect 560394 346054 561014 381498
rect 560394 345498 560426 346054
rect 560982 345498 561014 346054
rect 560394 310054 561014 345498
rect 560394 309498 560426 310054
rect 560982 309498 561014 310054
rect 560394 274054 561014 309498
rect 560394 273498 560426 274054
rect 560982 273498 561014 274054
rect 560394 238054 561014 273498
rect 560394 237498 560426 238054
rect 560982 237498 561014 238054
rect 560394 202054 561014 237498
rect 560394 201498 560426 202054
rect 560982 201498 561014 202054
rect 560394 166054 561014 201498
rect 560394 165498 560426 166054
rect 560982 165498 561014 166054
rect 560394 130054 561014 165498
rect 560394 129498 560426 130054
rect 560982 129498 561014 130054
rect 560394 94054 561014 129498
rect 560394 93498 560426 94054
rect 560982 93498 561014 94054
rect 560394 58054 561014 93498
rect 560394 57498 560426 58054
rect 560982 57498 561014 58054
rect 560394 22054 561014 57498
rect 560394 21498 560426 22054
rect 560982 21498 561014 22054
rect 560394 -5146 561014 21498
rect 560394 -5702 560426 -5146
rect 560982 -5702 561014 -5146
rect 560394 -7654 561014 -5702
rect 564114 710598 564734 711590
rect 564114 710042 564146 710598
rect 564702 710042 564734 710598
rect 564114 673774 564734 710042
rect 564114 673218 564146 673774
rect 564702 673218 564734 673774
rect 564114 637774 564734 673218
rect 564114 637218 564146 637774
rect 564702 637218 564734 637774
rect 564114 601774 564734 637218
rect 564114 601218 564146 601774
rect 564702 601218 564734 601774
rect 564114 565774 564734 601218
rect 564114 565218 564146 565774
rect 564702 565218 564734 565774
rect 564114 529774 564734 565218
rect 564114 529218 564146 529774
rect 564702 529218 564734 529774
rect 564114 493774 564734 529218
rect 564114 493218 564146 493774
rect 564702 493218 564734 493774
rect 564114 457774 564734 493218
rect 564114 457218 564146 457774
rect 564702 457218 564734 457774
rect 564114 421774 564734 457218
rect 564114 421218 564146 421774
rect 564702 421218 564734 421774
rect 564114 385774 564734 421218
rect 564114 385218 564146 385774
rect 564702 385218 564734 385774
rect 564114 349774 564734 385218
rect 564114 349218 564146 349774
rect 564702 349218 564734 349774
rect 564114 313774 564734 349218
rect 564114 313218 564146 313774
rect 564702 313218 564734 313774
rect 564114 277774 564734 313218
rect 564114 277218 564146 277774
rect 564702 277218 564734 277774
rect 564114 241774 564734 277218
rect 564114 241218 564146 241774
rect 564702 241218 564734 241774
rect 564114 205774 564734 241218
rect 564114 205218 564146 205774
rect 564702 205218 564734 205774
rect 564114 169774 564734 205218
rect 564114 169218 564146 169774
rect 564702 169218 564734 169774
rect 564114 133774 564734 169218
rect 564114 133218 564146 133774
rect 564702 133218 564734 133774
rect 564114 97774 564734 133218
rect 564114 97218 564146 97774
rect 564702 97218 564734 97774
rect 564114 61774 564734 97218
rect 564114 61218 564146 61774
rect 564702 61218 564734 61774
rect 564114 25774 564734 61218
rect 564114 25218 564146 25774
rect 564702 25218 564734 25774
rect 564114 -6106 564734 25218
rect 564114 -6662 564146 -6106
rect 564702 -6662 564734 -6106
rect 564114 -7654 564734 -6662
rect 567834 711558 568454 711590
rect 567834 711002 567866 711558
rect 568422 711002 568454 711558
rect 567834 677494 568454 711002
rect 567834 676938 567866 677494
rect 568422 676938 568454 677494
rect 567834 641494 568454 676938
rect 567834 640938 567866 641494
rect 568422 640938 568454 641494
rect 567834 605494 568454 640938
rect 567834 604938 567866 605494
rect 568422 604938 568454 605494
rect 567834 569494 568454 604938
rect 567834 568938 567866 569494
rect 568422 568938 568454 569494
rect 567834 533494 568454 568938
rect 567834 532938 567866 533494
rect 568422 532938 568454 533494
rect 567834 497494 568454 532938
rect 567834 496938 567866 497494
rect 568422 496938 568454 497494
rect 567834 461494 568454 496938
rect 567834 460938 567866 461494
rect 568422 460938 568454 461494
rect 567834 425494 568454 460938
rect 567834 424938 567866 425494
rect 568422 424938 568454 425494
rect 567834 389494 568454 424938
rect 567834 388938 567866 389494
rect 568422 388938 568454 389494
rect 567834 353494 568454 388938
rect 567834 352938 567866 353494
rect 568422 352938 568454 353494
rect 567834 317494 568454 352938
rect 577794 704838 578414 711590
rect 577794 704282 577826 704838
rect 578382 704282 578414 704838
rect 577794 687454 578414 704282
rect 577794 686898 577826 687454
rect 578382 686898 578414 687454
rect 577794 651454 578414 686898
rect 577794 650898 577826 651454
rect 578382 650898 578414 651454
rect 577794 615454 578414 650898
rect 577794 614898 577826 615454
rect 578382 614898 578414 615454
rect 577794 579454 578414 614898
rect 577794 578898 577826 579454
rect 578382 578898 578414 579454
rect 577794 543454 578414 578898
rect 577794 542898 577826 543454
rect 578382 542898 578414 543454
rect 577794 507454 578414 542898
rect 577794 506898 577826 507454
rect 578382 506898 578414 507454
rect 577794 471454 578414 506898
rect 577794 470898 577826 471454
rect 578382 470898 578414 471454
rect 577794 435454 578414 470898
rect 577794 434898 577826 435454
rect 578382 434898 578414 435454
rect 577794 399454 578414 434898
rect 577794 398898 577826 399454
rect 578382 398898 578414 399454
rect 577794 363454 578414 398898
rect 577794 362898 577826 363454
rect 578382 362898 578414 363454
rect 569168 327454 569488 327486
rect 569168 327218 569210 327454
rect 569446 327218 569488 327454
rect 569168 327134 569488 327218
rect 569168 326898 569210 327134
rect 569446 326898 569488 327134
rect 569168 326866 569488 326898
rect 577794 327454 578414 362898
rect 577794 326898 577826 327454
rect 578382 326898 578414 327454
rect 567834 316938 567866 317494
rect 568422 316938 568454 317494
rect 567834 281494 568454 316938
rect 569168 291454 569488 291486
rect 569168 291218 569210 291454
rect 569446 291218 569488 291454
rect 569168 291134 569488 291218
rect 569168 290898 569210 291134
rect 569446 290898 569488 291134
rect 569168 290866 569488 290898
rect 577794 291454 578414 326898
rect 577794 290898 577826 291454
rect 578382 290898 578414 291454
rect 567834 280938 567866 281494
rect 568422 280938 568454 281494
rect 567834 245494 568454 280938
rect 569168 255454 569488 255486
rect 569168 255218 569210 255454
rect 569446 255218 569488 255454
rect 569168 255134 569488 255218
rect 569168 254898 569210 255134
rect 569446 254898 569488 255134
rect 569168 254866 569488 254898
rect 577794 255454 578414 290898
rect 577794 254898 577826 255454
rect 578382 254898 578414 255454
rect 567834 244938 567866 245494
rect 568422 244938 568454 245494
rect 567834 209494 568454 244938
rect 569168 219454 569488 219486
rect 569168 219218 569210 219454
rect 569446 219218 569488 219454
rect 569168 219134 569488 219218
rect 569168 218898 569210 219134
rect 569446 218898 569488 219134
rect 569168 218866 569488 218898
rect 577794 219454 578414 254898
rect 577794 218898 577826 219454
rect 578382 218898 578414 219454
rect 567834 208938 567866 209494
rect 568422 208938 568454 209494
rect 567834 173494 568454 208938
rect 569168 183454 569488 183486
rect 569168 183218 569210 183454
rect 569446 183218 569488 183454
rect 569168 183134 569488 183218
rect 569168 182898 569210 183134
rect 569446 182898 569488 183134
rect 569168 182866 569488 182898
rect 577794 183454 578414 218898
rect 577794 182898 577826 183454
rect 578382 182898 578414 183454
rect 567834 172938 567866 173494
rect 568422 172938 568454 173494
rect 567834 137494 568454 172938
rect 569168 147454 569488 147486
rect 569168 147218 569210 147454
rect 569446 147218 569488 147454
rect 569168 147134 569488 147218
rect 569168 146898 569210 147134
rect 569446 146898 569488 147134
rect 569168 146866 569488 146898
rect 577794 147454 578414 182898
rect 577794 146898 577826 147454
rect 578382 146898 578414 147454
rect 567834 136938 567866 137494
rect 568422 136938 568454 137494
rect 567834 101494 568454 136938
rect 569168 111454 569488 111486
rect 569168 111218 569210 111454
rect 569446 111218 569488 111454
rect 569168 111134 569488 111218
rect 569168 110898 569210 111134
rect 569446 110898 569488 111134
rect 569168 110866 569488 110898
rect 577794 111454 578414 146898
rect 577794 110898 577826 111454
rect 578382 110898 578414 111454
rect 567834 100938 567866 101494
rect 568422 100938 568454 101494
rect 567834 65494 568454 100938
rect 569168 75454 569488 75486
rect 569168 75218 569210 75454
rect 569446 75218 569488 75454
rect 569168 75134 569488 75218
rect 569168 74898 569210 75134
rect 569446 74898 569488 75134
rect 569168 74866 569488 74898
rect 577794 75454 578414 110898
rect 577794 74898 577826 75454
rect 578382 74898 578414 75454
rect 567834 64938 567866 65494
rect 568422 64938 568454 65494
rect 567834 29494 568454 64938
rect 569168 39454 569488 39486
rect 569168 39218 569210 39454
rect 569446 39218 569488 39454
rect 569168 39134 569488 39218
rect 569168 38898 569210 39134
rect 569446 38898 569488 39134
rect 569168 38866 569488 38898
rect 577794 39454 578414 74898
rect 577794 38898 577826 39454
rect 578382 38898 578414 39454
rect 567834 28938 567866 29494
rect 568422 28938 568454 29494
rect 567834 -7066 568454 28938
rect 567834 -7622 567866 -7066
rect 568422 -7622 568454 -7066
rect 567834 -7654 568454 -7622
rect 577794 3454 578414 38898
rect 577794 2898 577826 3454
rect 578382 2898 578414 3454
rect 577794 -346 578414 2898
rect 577794 -902 577826 -346
rect 578382 -902 578414 -346
rect 577794 -7654 578414 -902
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711002 592062 711558
rect 592618 711002 592650 711558
rect 591070 710598 591690 710630
rect 591070 710042 591102 710598
rect 591658 710042 591690 710598
rect 590110 709638 590730 709670
rect 590110 709082 590142 709638
rect 590698 709082 590730 709638
rect 589150 708678 589770 708710
rect 589150 708122 589182 708678
rect 589738 708122 589770 708678
rect 588190 707718 588810 707750
rect 588190 707162 588222 707718
rect 588778 707162 588810 707718
rect 587230 706758 587850 706790
rect 587230 706202 587262 706758
rect 587818 706202 587850 706758
rect 581514 705242 581546 705798
rect 582102 705242 582134 705798
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705242 586302 705798
rect 586858 705242 586890 705798
rect 581514 690618 581546 691174
rect 582102 690618 582134 691174
rect 581514 655174 582134 690618
rect 581514 654618 581546 655174
rect 582102 654618 582134 655174
rect 581514 619174 582134 654618
rect 581514 618618 581546 619174
rect 582102 618618 582134 619174
rect 581514 583174 582134 618618
rect 581514 582618 581546 583174
rect 582102 582618 582134 583174
rect 581514 547174 582134 582618
rect 581514 546618 581546 547174
rect 582102 546618 582134 547174
rect 581514 511174 582134 546618
rect 581514 510618 581546 511174
rect 582102 510618 582134 511174
rect 581514 475174 582134 510618
rect 581514 474618 581546 475174
rect 582102 474618 582134 475174
rect 581514 439174 582134 474618
rect 581514 438618 581546 439174
rect 582102 438618 582134 439174
rect 581514 403174 582134 438618
rect 581514 402618 581546 403174
rect 582102 402618 582134 403174
rect 581514 367174 582134 402618
rect 581514 366618 581546 367174
rect 582102 366618 582134 367174
rect 581514 331174 582134 366618
rect 581514 330618 581546 331174
rect 582102 330618 582134 331174
rect 581514 295174 582134 330618
rect 581514 294618 581546 295174
rect 582102 294618 582134 295174
rect 581514 259174 582134 294618
rect 581514 258618 581546 259174
rect 582102 258618 582134 259174
rect 581514 223174 582134 258618
rect 581514 222618 581546 223174
rect 582102 222618 582134 223174
rect 581514 187174 582134 222618
rect 581514 186618 581546 187174
rect 582102 186618 582134 187174
rect 581514 151174 582134 186618
rect 581514 150618 581546 151174
rect 582102 150618 582134 151174
rect 581514 115174 582134 150618
rect 581514 114618 581546 115174
rect 582102 114618 582134 115174
rect 581514 79174 582134 114618
rect 581514 78618 581546 79174
rect 582102 78618 582134 79174
rect 581514 43174 582134 78618
rect 581514 42618 581546 43174
rect 582102 42618 582134 43174
rect 581514 7174 582134 42618
rect 581514 6618 581546 7174
rect 582102 6618 582134 7174
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704282 585342 704838
rect 585898 704282 585930 704838
rect 585310 687454 585930 704282
rect 585310 686898 585342 687454
rect 585898 686898 585930 687454
rect 585310 651454 585930 686898
rect 585310 650898 585342 651454
rect 585898 650898 585930 651454
rect 585310 615454 585930 650898
rect 585310 614898 585342 615454
rect 585898 614898 585930 615454
rect 585310 579454 585930 614898
rect 585310 578898 585342 579454
rect 585898 578898 585930 579454
rect 585310 543454 585930 578898
rect 585310 542898 585342 543454
rect 585898 542898 585930 543454
rect 585310 507454 585930 542898
rect 585310 506898 585342 507454
rect 585898 506898 585930 507454
rect 585310 471454 585930 506898
rect 585310 470898 585342 471454
rect 585898 470898 585930 471454
rect 585310 435454 585930 470898
rect 585310 434898 585342 435454
rect 585898 434898 585930 435454
rect 585310 399454 585930 434898
rect 585310 398898 585342 399454
rect 585898 398898 585930 399454
rect 585310 363454 585930 398898
rect 585310 362898 585342 363454
rect 585898 362898 585930 363454
rect 585310 327454 585930 362898
rect 585310 326898 585342 327454
rect 585898 326898 585930 327454
rect 585310 291454 585930 326898
rect 585310 290898 585342 291454
rect 585898 290898 585930 291454
rect 585310 255454 585930 290898
rect 585310 254898 585342 255454
rect 585898 254898 585930 255454
rect 585310 219454 585930 254898
rect 585310 218898 585342 219454
rect 585898 218898 585930 219454
rect 585310 183454 585930 218898
rect 585310 182898 585342 183454
rect 585898 182898 585930 183454
rect 585310 147454 585930 182898
rect 585310 146898 585342 147454
rect 585898 146898 585930 147454
rect 585310 111454 585930 146898
rect 585310 110898 585342 111454
rect 585898 110898 585930 111454
rect 585310 75454 585930 110898
rect 585310 74898 585342 75454
rect 585898 74898 585930 75454
rect 585310 39454 585930 74898
rect 585310 38898 585342 39454
rect 585898 38898 585930 39454
rect 585310 3454 585930 38898
rect 585310 2898 585342 3454
rect 585898 2898 585930 3454
rect 585310 -346 585930 2898
rect 585310 -902 585342 -346
rect 585898 -902 585930 -346
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690618 586302 691174
rect 586858 690618 586890 691174
rect 586270 655174 586890 690618
rect 586270 654618 586302 655174
rect 586858 654618 586890 655174
rect 586270 619174 586890 654618
rect 586270 618618 586302 619174
rect 586858 618618 586890 619174
rect 586270 583174 586890 618618
rect 586270 582618 586302 583174
rect 586858 582618 586890 583174
rect 586270 547174 586890 582618
rect 586270 546618 586302 547174
rect 586858 546618 586890 547174
rect 586270 511174 586890 546618
rect 586270 510618 586302 511174
rect 586858 510618 586890 511174
rect 586270 475174 586890 510618
rect 586270 474618 586302 475174
rect 586858 474618 586890 475174
rect 586270 439174 586890 474618
rect 586270 438618 586302 439174
rect 586858 438618 586890 439174
rect 586270 403174 586890 438618
rect 586270 402618 586302 403174
rect 586858 402618 586890 403174
rect 586270 367174 586890 402618
rect 586270 366618 586302 367174
rect 586858 366618 586890 367174
rect 586270 331174 586890 366618
rect 586270 330618 586302 331174
rect 586858 330618 586890 331174
rect 586270 295174 586890 330618
rect 586270 294618 586302 295174
rect 586858 294618 586890 295174
rect 586270 259174 586890 294618
rect 586270 258618 586302 259174
rect 586858 258618 586890 259174
rect 586270 223174 586890 258618
rect 586270 222618 586302 223174
rect 586858 222618 586890 223174
rect 586270 187174 586890 222618
rect 586270 186618 586302 187174
rect 586858 186618 586890 187174
rect 586270 151174 586890 186618
rect 586270 150618 586302 151174
rect 586858 150618 586890 151174
rect 586270 115174 586890 150618
rect 586270 114618 586302 115174
rect 586858 114618 586890 115174
rect 586270 79174 586890 114618
rect 586270 78618 586302 79174
rect 586858 78618 586890 79174
rect 586270 43174 586890 78618
rect 586270 42618 586302 43174
rect 586858 42618 586890 43174
rect 586270 7174 586890 42618
rect 586270 6618 586302 7174
rect 586858 6618 586890 7174
rect 581514 -1862 581546 -1306
rect 582102 -1862 582134 -1306
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1862 586302 -1306
rect 586858 -1862 586890 -1306
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694338 587262 694894
rect 587818 694338 587850 694894
rect 587230 658894 587850 694338
rect 587230 658338 587262 658894
rect 587818 658338 587850 658894
rect 587230 622894 587850 658338
rect 587230 622338 587262 622894
rect 587818 622338 587850 622894
rect 587230 586894 587850 622338
rect 587230 586338 587262 586894
rect 587818 586338 587850 586894
rect 587230 550894 587850 586338
rect 587230 550338 587262 550894
rect 587818 550338 587850 550894
rect 587230 514894 587850 550338
rect 587230 514338 587262 514894
rect 587818 514338 587850 514894
rect 587230 478894 587850 514338
rect 587230 478338 587262 478894
rect 587818 478338 587850 478894
rect 587230 442894 587850 478338
rect 587230 442338 587262 442894
rect 587818 442338 587850 442894
rect 587230 406894 587850 442338
rect 587230 406338 587262 406894
rect 587818 406338 587850 406894
rect 587230 370894 587850 406338
rect 587230 370338 587262 370894
rect 587818 370338 587850 370894
rect 587230 334894 587850 370338
rect 587230 334338 587262 334894
rect 587818 334338 587850 334894
rect 587230 298894 587850 334338
rect 587230 298338 587262 298894
rect 587818 298338 587850 298894
rect 587230 262894 587850 298338
rect 587230 262338 587262 262894
rect 587818 262338 587850 262894
rect 587230 226894 587850 262338
rect 587230 226338 587262 226894
rect 587818 226338 587850 226894
rect 587230 190894 587850 226338
rect 587230 190338 587262 190894
rect 587818 190338 587850 190894
rect 587230 154894 587850 190338
rect 587230 154338 587262 154894
rect 587818 154338 587850 154894
rect 587230 118894 587850 154338
rect 587230 118338 587262 118894
rect 587818 118338 587850 118894
rect 587230 82894 587850 118338
rect 587230 82338 587262 82894
rect 587818 82338 587850 82894
rect 587230 46894 587850 82338
rect 587230 46338 587262 46894
rect 587818 46338 587850 46894
rect 587230 10894 587850 46338
rect 587230 10338 587262 10894
rect 587818 10338 587850 10894
rect 587230 -2266 587850 10338
rect 587230 -2822 587262 -2266
rect 587818 -2822 587850 -2266
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698058 588222 698614
rect 588778 698058 588810 698614
rect 588190 662614 588810 698058
rect 588190 662058 588222 662614
rect 588778 662058 588810 662614
rect 588190 626614 588810 662058
rect 588190 626058 588222 626614
rect 588778 626058 588810 626614
rect 588190 590614 588810 626058
rect 588190 590058 588222 590614
rect 588778 590058 588810 590614
rect 588190 554614 588810 590058
rect 588190 554058 588222 554614
rect 588778 554058 588810 554614
rect 588190 518614 588810 554058
rect 588190 518058 588222 518614
rect 588778 518058 588810 518614
rect 588190 482614 588810 518058
rect 588190 482058 588222 482614
rect 588778 482058 588810 482614
rect 588190 446614 588810 482058
rect 588190 446058 588222 446614
rect 588778 446058 588810 446614
rect 588190 410614 588810 446058
rect 588190 410058 588222 410614
rect 588778 410058 588810 410614
rect 588190 374614 588810 410058
rect 588190 374058 588222 374614
rect 588778 374058 588810 374614
rect 588190 338614 588810 374058
rect 588190 338058 588222 338614
rect 588778 338058 588810 338614
rect 588190 302614 588810 338058
rect 588190 302058 588222 302614
rect 588778 302058 588810 302614
rect 588190 266614 588810 302058
rect 588190 266058 588222 266614
rect 588778 266058 588810 266614
rect 588190 230614 588810 266058
rect 588190 230058 588222 230614
rect 588778 230058 588810 230614
rect 588190 194614 588810 230058
rect 588190 194058 588222 194614
rect 588778 194058 588810 194614
rect 588190 158614 588810 194058
rect 588190 158058 588222 158614
rect 588778 158058 588810 158614
rect 588190 122614 588810 158058
rect 588190 122058 588222 122614
rect 588778 122058 588810 122614
rect 588190 86614 588810 122058
rect 588190 86058 588222 86614
rect 588778 86058 588810 86614
rect 588190 50614 588810 86058
rect 588190 50058 588222 50614
rect 588778 50058 588810 50614
rect 588190 14614 588810 50058
rect 588190 14058 588222 14614
rect 588778 14058 588810 14614
rect 588190 -3226 588810 14058
rect 588190 -3782 588222 -3226
rect 588778 -3782 588810 -3226
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 665778 589182 666334
rect 589738 665778 589770 666334
rect 589150 630334 589770 665778
rect 589150 629778 589182 630334
rect 589738 629778 589770 630334
rect 589150 594334 589770 629778
rect 589150 593778 589182 594334
rect 589738 593778 589770 594334
rect 589150 558334 589770 593778
rect 589150 557778 589182 558334
rect 589738 557778 589770 558334
rect 589150 522334 589770 557778
rect 589150 521778 589182 522334
rect 589738 521778 589770 522334
rect 589150 486334 589770 521778
rect 589150 485778 589182 486334
rect 589738 485778 589770 486334
rect 589150 450334 589770 485778
rect 589150 449778 589182 450334
rect 589738 449778 589770 450334
rect 589150 414334 589770 449778
rect 589150 413778 589182 414334
rect 589738 413778 589770 414334
rect 589150 378334 589770 413778
rect 589150 377778 589182 378334
rect 589738 377778 589770 378334
rect 589150 342334 589770 377778
rect 589150 341778 589182 342334
rect 589738 341778 589770 342334
rect 589150 306334 589770 341778
rect 589150 305778 589182 306334
rect 589738 305778 589770 306334
rect 589150 270334 589770 305778
rect 589150 269778 589182 270334
rect 589738 269778 589770 270334
rect 589150 234334 589770 269778
rect 589150 233778 589182 234334
rect 589738 233778 589770 234334
rect 589150 198334 589770 233778
rect 589150 197778 589182 198334
rect 589738 197778 589770 198334
rect 589150 162334 589770 197778
rect 589150 161778 589182 162334
rect 589738 161778 589770 162334
rect 589150 126334 589770 161778
rect 589150 125778 589182 126334
rect 589738 125778 589770 126334
rect 589150 90334 589770 125778
rect 589150 89778 589182 90334
rect 589738 89778 589770 90334
rect 589150 54334 589770 89778
rect 589150 53778 589182 54334
rect 589738 53778 589770 54334
rect 589150 18334 589770 53778
rect 589150 17778 589182 18334
rect 589738 17778 589770 18334
rect 589150 -4186 589770 17778
rect 589150 -4742 589182 -4186
rect 589738 -4742 589770 -4186
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669498 590142 670054
rect 590698 669498 590730 670054
rect 590110 634054 590730 669498
rect 590110 633498 590142 634054
rect 590698 633498 590730 634054
rect 590110 598054 590730 633498
rect 590110 597498 590142 598054
rect 590698 597498 590730 598054
rect 590110 562054 590730 597498
rect 590110 561498 590142 562054
rect 590698 561498 590730 562054
rect 590110 526054 590730 561498
rect 590110 525498 590142 526054
rect 590698 525498 590730 526054
rect 590110 490054 590730 525498
rect 590110 489498 590142 490054
rect 590698 489498 590730 490054
rect 590110 454054 590730 489498
rect 590110 453498 590142 454054
rect 590698 453498 590730 454054
rect 590110 418054 590730 453498
rect 590110 417498 590142 418054
rect 590698 417498 590730 418054
rect 590110 382054 590730 417498
rect 590110 381498 590142 382054
rect 590698 381498 590730 382054
rect 590110 346054 590730 381498
rect 590110 345498 590142 346054
rect 590698 345498 590730 346054
rect 590110 310054 590730 345498
rect 590110 309498 590142 310054
rect 590698 309498 590730 310054
rect 590110 274054 590730 309498
rect 590110 273498 590142 274054
rect 590698 273498 590730 274054
rect 590110 238054 590730 273498
rect 590110 237498 590142 238054
rect 590698 237498 590730 238054
rect 590110 202054 590730 237498
rect 590110 201498 590142 202054
rect 590698 201498 590730 202054
rect 590110 166054 590730 201498
rect 590110 165498 590142 166054
rect 590698 165498 590730 166054
rect 590110 130054 590730 165498
rect 590110 129498 590142 130054
rect 590698 129498 590730 130054
rect 590110 94054 590730 129498
rect 590110 93498 590142 94054
rect 590698 93498 590730 94054
rect 590110 58054 590730 93498
rect 590110 57498 590142 58054
rect 590698 57498 590730 58054
rect 590110 22054 590730 57498
rect 590110 21498 590142 22054
rect 590698 21498 590730 22054
rect 590110 -5146 590730 21498
rect 590110 -5702 590142 -5146
rect 590698 -5702 590730 -5146
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673218 591102 673774
rect 591658 673218 591690 673774
rect 591070 637774 591690 673218
rect 591070 637218 591102 637774
rect 591658 637218 591690 637774
rect 591070 601774 591690 637218
rect 591070 601218 591102 601774
rect 591658 601218 591690 601774
rect 591070 565774 591690 601218
rect 591070 565218 591102 565774
rect 591658 565218 591690 565774
rect 591070 529774 591690 565218
rect 591070 529218 591102 529774
rect 591658 529218 591690 529774
rect 591070 493774 591690 529218
rect 591070 493218 591102 493774
rect 591658 493218 591690 493774
rect 591070 457774 591690 493218
rect 591070 457218 591102 457774
rect 591658 457218 591690 457774
rect 591070 421774 591690 457218
rect 591070 421218 591102 421774
rect 591658 421218 591690 421774
rect 591070 385774 591690 421218
rect 591070 385218 591102 385774
rect 591658 385218 591690 385774
rect 591070 349774 591690 385218
rect 591070 349218 591102 349774
rect 591658 349218 591690 349774
rect 591070 313774 591690 349218
rect 591070 313218 591102 313774
rect 591658 313218 591690 313774
rect 591070 277774 591690 313218
rect 591070 277218 591102 277774
rect 591658 277218 591690 277774
rect 591070 241774 591690 277218
rect 591070 241218 591102 241774
rect 591658 241218 591690 241774
rect 591070 205774 591690 241218
rect 591070 205218 591102 205774
rect 591658 205218 591690 205774
rect 591070 169774 591690 205218
rect 591070 169218 591102 169774
rect 591658 169218 591690 169774
rect 591070 133774 591690 169218
rect 591070 133218 591102 133774
rect 591658 133218 591690 133774
rect 591070 97774 591690 133218
rect 591070 97218 591102 97774
rect 591658 97218 591690 97774
rect 591070 61774 591690 97218
rect 591070 61218 591102 61774
rect 591658 61218 591690 61774
rect 591070 25774 591690 61218
rect 591070 25218 591102 25774
rect 591658 25218 591690 25774
rect 591070 -6106 591690 25218
rect 591070 -6662 591102 -6106
rect 591658 -6662 591690 -6106
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 676938 592062 677494
rect 592618 676938 592650 677494
rect 592030 641494 592650 676938
rect 592030 640938 592062 641494
rect 592618 640938 592650 641494
rect 592030 605494 592650 640938
rect 592030 604938 592062 605494
rect 592618 604938 592650 605494
rect 592030 569494 592650 604938
rect 592030 568938 592062 569494
rect 592618 568938 592650 569494
rect 592030 533494 592650 568938
rect 592030 532938 592062 533494
rect 592618 532938 592650 533494
rect 592030 497494 592650 532938
rect 592030 496938 592062 497494
rect 592618 496938 592650 497494
rect 592030 461494 592650 496938
rect 592030 460938 592062 461494
rect 592618 460938 592650 461494
rect 592030 425494 592650 460938
rect 592030 424938 592062 425494
rect 592618 424938 592650 425494
rect 592030 389494 592650 424938
rect 592030 388938 592062 389494
rect 592618 388938 592650 389494
rect 592030 353494 592650 388938
rect 592030 352938 592062 353494
rect 592618 352938 592650 353494
rect 592030 317494 592650 352938
rect 592030 316938 592062 317494
rect 592618 316938 592650 317494
rect 592030 281494 592650 316938
rect 592030 280938 592062 281494
rect 592618 280938 592650 281494
rect 592030 245494 592650 280938
rect 592030 244938 592062 245494
rect 592618 244938 592650 245494
rect 592030 209494 592650 244938
rect 592030 208938 592062 209494
rect 592618 208938 592650 209494
rect 592030 173494 592650 208938
rect 592030 172938 592062 173494
rect 592618 172938 592650 173494
rect 592030 137494 592650 172938
rect 592030 136938 592062 137494
rect 592618 136938 592650 137494
rect 592030 101494 592650 136938
rect 592030 100938 592062 101494
rect 592618 100938 592650 101494
rect 592030 65494 592650 100938
rect 592030 64938 592062 65494
rect 592618 64938 592650 65494
rect 592030 29494 592650 64938
rect 592030 28938 592062 29494
rect 592618 28938 592650 29494
rect 592030 -7066 592650 28938
rect 592030 -7622 592062 -7066
rect 592618 -7622 592650 -7066
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711002 -8138 711558
rect -8694 676938 -8138 677494
rect -8694 640938 -8138 641494
rect -8694 604938 -8138 605494
rect -8694 568938 -8138 569494
rect -8694 532938 -8138 533494
rect -8694 496938 -8138 497494
rect -8694 460938 -8138 461494
rect -8694 424938 -8138 425494
rect -8694 388938 -8138 389494
rect -8694 352938 -8138 353494
rect -8694 316938 -8138 317494
rect -8694 280938 -8138 281494
rect -8694 244938 -8138 245494
rect -8694 208938 -8138 209494
rect -8694 172938 -8138 173494
rect -8694 136938 -8138 137494
rect -8694 100938 -8138 101494
rect -8694 64938 -8138 65494
rect -8694 28938 -8138 29494
rect -7734 710042 -7178 710598
rect -7734 673218 -7178 673774
rect -7734 637218 -7178 637774
rect -7734 601218 -7178 601774
rect -7734 565218 -7178 565774
rect -7734 529218 -7178 529774
rect -7734 493218 -7178 493774
rect -7734 457218 -7178 457774
rect -7734 421218 -7178 421774
rect -7734 385218 -7178 385774
rect -7734 349218 -7178 349774
rect -7734 313218 -7178 313774
rect -7734 277218 -7178 277774
rect -7734 241218 -7178 241774
rect -7734 205218 -7178 205774
rect -7734 169218 -7178 169774
rect -7734 133218 -7178 133774
rect -7734 97218 -7178 97774
rect -7734 61218 -7178 61774
rect -7734 25218 -7178 25774
rect -6774 709082 -6218 709638
rect -6774 669498 -6218 670054
rect -6774 633498 -6218 634054
rect -6774 597498 -6218 598054
rect -6774 561498 -6218 562054
rect -6774 525498 -6218 526054
rect -6774 489498 -6218 490054
rect -6774 453498 -6218 454054
rect -6774 417498 -6218 418054
rect -6774 381498 -6218 382054
rect -6774 345498 -6218 346054
rect -6774 309498 -6218 310054
rect -6774 273498 -6218 274054
rect -6774 237498 -6218 238054
rect -6774 201498 -6218 202054
rect -6774 165498 -6218 166054
rect -6774 129498 -6218 130054
rect -6774 93498 -6218 94054
rect -6774 57498 -6218 58054
rect -6774 21498 -6218 22054
rect -5814 708122 -5258 708678
rect -5814 665778 -5258 666334
rect -5814 629778 -5258 630334
rect -5814 593778 -5258 594334
rect -5814 557778 -5258 558334
rect -5814 521778 -5258 522334
rect -5814 485778 -5258 486334
rect -5814 449778 -5258 450334
rect -5814 413778 -5258 414334
rect -5814 377778 -5258 378334
rect -5814 341778 -5258 342334
rect -5814 305778 -5258 306334
rect -5814 269778 -5258 270334
rect -5814 233778 -5258 234334
rect -5814 197778 -5258 198334
rect -5814 161778 -5258 162334
rect -5814 125778 -5258 126334
rect -5814 89778 -5258 90334
rect -5814 53778 -5258 54334
rect -5814 17778 -5258 18334
rect -4854 707162 -4298 707718
rect -4854 698058 -4298 698614
rect -4854 662058 -4298 662614
rect -4854 626058 -4298 626614
rect -4854 590058 -4298 590614
rect -4854 554058 -4298 554614
rect -4854 518058 -4298 518614
rect -4854 482058 -4298 482614
rect -4854 446058 -4298 446614
rect -4854 410058 -4298 410614
rect -4854 374058 -4298 374614
rect -4854 338058 -4298 338614
rect -4854 302058 -4298 302614
rect -4854 266058 -4298 266614
rect -4854 230058 -4298 230614
rect -4854 194058 -4298 194614
rect -4854 158058 -4298 158614
rect -4854 122058 -4298 122614
rect -4854 86058 -4298 86614
rect -4854 50058 -4298 50614
rect -4854 14058 -4298 14614
rect -3894 706202 -3338 706758
rect -3894 694338 -3338 694894
rect -3894 658338 -3338 658894
rect -3894 622338 -3338 622894
rect -3894 586338 -3338 586894
rect -3894 550338 -3338 550894
rect -3894 514338 -3338 514894
rect -3894 478338 -3338 478894
rect -3894 442338 -3338 442894
rect -3894 406338 -3338 406894
rect -3894 370338 -3338 370894
rect -3894 334338 -3338 334894
rect -3894 298338 -3338 298894
rect -3894 262338 -3338 262894
rect -3894 226338 -3338 226894
rect -3894 190338 -3338 190894
rect -3894 154338 -3338 154894
rect -3894 118338 -3338 118894
rect -3894 82338 -3338 82894
rect -3894 46338 -3338 46894
rect -3894 10338 -3338 10894
rect -2934 705242 -2378 705798
rect -2934 690618 -2378 691174
rect -2934 654618 -2378 655174
rect -2934 618618 -2378 619174
rect -2934 582618 -2378 583174
rect -2934 546618 -2378 547174
rect -2934 510618 -2378 511174
rect -2934 474618 -2378 475174
rect -2934 438618 -2378 439174
rect -2934 402618 -2378 403174
rect -2934 366618 -2378 367174
rect -2934 330618 -2378 331174
rect -2934 294618 -2378 295174
rect -2934 258618 -2378 259174
rect -2934 222618 -2378 223174
rect -2934 186618 -2378 187174
rect -2934 150618 -2378 151174
rect -2934 114618 -2378 115174
rect -2934 78618 -2378 79174
rect -2934 42618 -2378 43174
rect -2934 6618 -2378 7174
rect -1974 704282 -1418 704838
rect -1974 686898 -1418 687454
rect -1974 650898 -1418 651454
rect -1974 614898 -1418 615454
rect -1974 578898 -1418 579454
rect -1974 542898 -1418 543454
rect -1974 506898 -1418 507454
rect -1974 470898 -1418 471454
rect -1974 434898 -1418 435454
rect -1974 398898 -1418 399454
rect -1974 362898 -1418 363454
rect -1974 326898 -1418 327454
rect -1974 290898 -1418 291454
rect -1974 254898 -1418 255454
rect -1974 218898 -1418 219454
rect -1974 182898 -1418 183454
rect -1974 146898 -1418 147454
rect -1974 110898 -1418 111454
rect -1974 74898 -1418 75454
rect -1974 38898 -1418 39454
rect -1974 2898 -1418 3454
rect -1974 -902 -1418 -346
rect 1826 704282 2382 704838
rect 1826 686898 2382 687454
rect 1826 650898 2382 651454
rect 1826 614898 2382 615454
rect 1826 578898 2382 579454
rect 1826 542898 2382 543454
rect 1826 506898 2382 507454
rect 1826 470898 2382 471454
rect 1826 434898 2382 435454
rect 1826 398898 2382 399454
rect 1826 362898 2382 363454
rect 1826 326898 2382 327454
rect 1826 290898 2382 291454
rect 1826 254898 2382 255454
rect 1826 218898 2382 219454
rect 1826 182898 2382 183454
rect 1826 146898 2382 147454
rect 1826 110898 2382 111454
rect 1826 74898 2382 75454
rect 1826 38898 2382 39454
rect 1826 2898 2382 3454
rect 1826 -902 2382 -346
rect -2934 -1862 -2378 -1306
rect -3894 -2822 -3338 -2266
rect -4854 -3782 -4298 -3226
rect -5814 -4742 -5258 -4186
rect -6774 -5702 -6218 -5146
rect -7734 -6662 -7178 -6106
rect -8694 -7622 -8138 -7066
rect 5546 705242 6102 705798
rect 5546 690618 6102 691174
rect 5546 654618 6102 655174
rect 5546 618618 6102 619174
rect 5546 582618 6102 583174
rect 5546 546618 6102 547174
rect 5546 510618 6102 511174
rect 5546 474618 6102 475174
rect 5546 438618 6102 439174
rect 5546 402618 6102 403174
rect 5546 366618 6102 367174
rect 5546 330618 6102 331174
rect 5546 294618 6102 295174
rect 5546 258618 6102 259174
rect 5546 222618 6102 223174
rect 5546 186618 6102 187174
rect 5546 150618 6102 151174
rect 5546 114618 6102 115174
rect 5546 78618 6102 79174
rect 5546 42618 6102 43174
rect 5546 6618 6102 7174
rect 5546 -1862 6102 -1306
rect 9266 706202 9822 706758
rect 9266 694338 9822 694894
rect 9266 658338 9822 658894
rect 9266 622338 9822 622894
rect 9266 586338 9822 586894
rect 9266 550338 9822 550894
rect 9266 514338 9822 514894
rect 9266 478338 9822 478894
rect 9266 442338 9822 442894
rect 9266 406338 9822 406894
rect 9266 370338 9822 370894
rect 9266 334338 9822 334894
rect 9266 298338 9822 298894
rect 9266 262338 9822 262894
rect 9266 226338 9822 226894
rect 9266 190338 9822 190894
rect 9266 154338 9822 154894
rect 9266 118338 9822 118894
rect 9266 82338 9822 82894
rect 9266 46338 9822 46894
rect 9266 10338 9822 10894
rect 9266 -2822 9822 -2266
rect 12986 707162 13542 707718
rect 12986 698058 13542 698614
rect 12986 662058 13542 662614
rect 12986 626058 13542 626614
rect 12986 590058 13542 590614
rect 12986 554058 13542 554614
rect 12986 518058 13542 518614
rect 12986 482058 13542 482614
rect 12986 446058 13542 446614
rect 12986 410058 13542 410614
rect 12986 374058 13542 374614
rect 12986 338058 13542 338614
rect 16706 708122 17262 708678
rect 16706 665778 17262 666334
rect 16706 629778 17262 630334
rect 16706 593778 17262 594334
rect 16706 557778 17262 558334
rect 16706 521778 17262 522334
rect 16706 485778 17262 486334
rect 16706 449778 17262 450334
rect 16706 413778 17262 414334
rect 16706 377778 17262 378334
rect 16706 341778 17262 342334
rect 16250 327218 16486 327454
rect 16250 326898 16486 327134
rect 12986 302058 13542 302614
rect 16706 305778 17262 306334
rect 16250 291218 16486 291454
rect 16250 290898 16486 291134
rect 12986 266058 13542 266614
rect 16706 269778 17262 270334
rect 16250 255218 16486 255454
rect 16250 254898 16486 255134
rect 12986 230058 13542 230614
rect 16706 233778 17262 234334
rect 16250 219218 16486 219454
rect 16250 218898 16486 219134
rect 12986 194058 13542 194614
rect 16706 197778 17262 198334
rect 16250 183218 16486 183454
rect 16250 182898 16486 183134
rect 12986 158058 13542 158614
rect 16706 161778 17262 162334
rect 16250 147218 16486 147454
rect 16250 146898 16486 147134
rect 12986 122058 13542 122614
rect 16706 125778 17262 126334
rect 16250 111218 16486 111454
rect 16250 110898 16486 111134
rect 12986 86058 13542 86614
rect 16706 89778 17262 90334
rect 16250 75218 16486 75454
rect 16250 74898 16486 75134
rect 12986 50058 13542 50614
rect 16706 53778 17262 54334
rect 16250 39218 16486 39454
rect 16250 38898 16486 39134
rect 12986 14058 13542 14614
rect 12986 -3782 13542 -3226
rect 16706 17778 17262 18334
rect 16706 -4742 17262 -4186
rect 20426 709082 20982 709638
rect 20426 669498 20982 670054
rect 20426 633498 20982 634054
rect 20426 597498 20982 598054
rect 20426 561498 20982 562054
rect 20426 525498 20982 526054
rect 20426 489498 20982 490054
rect 20426 453498 20982 454054
rect 20426 417498 20982 418054
rect 20426 381498 20982 382054
rect 20426 345498 20982 346054
rect 20426 309498 20982 310054
rect 20426 273498 20982 274054
rect 20426 237498 20982 238054
rect 20426 201498 20982 202054
rect 20426 165498 20982 166054
rect 20426 129498 20982 130054
rect 20426 93498 20982 94054
rect 20426 57498 20982 58054
rect 20426 21498 20982 22054
rect 20426 -5702 20982 -5146
rect 24146 710042 24702 710598
rect 24146 673218 24702 673774
rect 24146 637218 24702 637774
rect 24146 601218 24702 601774
rect 24146 565218 24702 565774
rect 24146 529218 24702 529774
rect 24146 493218 24702 493774
rect 24146 457218 24702 457774
rect 24146 421218 24702 421774
rect 24146 385218 24702 385774
rect 24146 349218 24702 349774
rect 24146 313218 24702 313774
rect 24146 277218 24702 277774
rect 24146 241218 24702 241774
rect 24146 205218 24702 205774
rect 24146 169218 24702 169774
rect 24146 133218 24702 133774
rect 24146 97218 24702 97774
rect 24146 61218 24702 61774
rect 24146 25218 24702 25774
rect 24146 -6662 24702 -6106
rect 27866 711002 28422 711558
rect 27866 676938 28422 677494
rect 27866 640938 28422 641494
rect 27866 604938 28422 605494
rect 27866 568938 28422 569494
rect 27866 532938 28422 533494
rect 27866 496938 28422 497494
rect 27866 460938 28422 461494
rect 27866 424938 28422 425494
rect 27866 388938 28422 389494
rect 27866 352938 28422 353494
rect 37826 704282 38382 704838
rect 37826 686898 38382 687454
rect 37826 650898 38382 651454
rect 37826 614898 38382 615454
rect 37826 578898 38382 579454
rect 37826 542898 38382 543454
rect 37826 506898 38382 507454
rect 37826 470898 38382 471454
rect 37826 434898 38382 435454
rect 37826 398898 38382 399454
rect 37826 362898 38382 363454
rect 31610 330938 31846 331174
rect 31610 330618 31846 330854
rect 27866 316938 28422 317494
rect 37826 326898 38382 327454
rect 31610 294938 31846 295174
rect 31610 294618 31846 294854
rect 27866 280938 28422 281494
rect 37826 290898 38382 291454
rect 31610 258938 31846 259174
rect 31610 258618 31846 258854
rect 27866 244938 28422 245494
rect 37826 254898 38382 255454
rect 31610 222938 31846 223174
rect 31610 222618 31846 222854
rect 27866 208938 28422 209494
rect 37826 218898 38382 219454
rect 31610 186938 31846 187174
rect 31610 186618 31846 186854
rect 27866 172938 28422 173494
rect 37826 182898 38382 183454
rect 31610 150938 31846 151174
rect 31610 150618 31846 150854
rect 27866 136938 28422 137494
rect 37826 146898 38382 147454
rect 31610 114938 31846 115174
rect 31610 114618 31846 114854
rect 27866 100938 28422 101494
rect 37826 110898 38382 111454
rect 31610 78938 31846 79174
rect 31610 78618 31846 78854
rect 27866 64938 28422 65494
rect 37826 74898 38382 75454
rect 31610 42938 31846 43174
rect 31610 42618 31846 42854
rect 27866 28938 28422 29494
rect 37826 38898 38382 39454
rect 31610 6938 31846 7174
rect 31610 6618 31846 6854
rect 27866 -7622 28422 -7066
rect 37826 2898 38382 3454
rect 37826 -902 38382 -346
rect 41546 705242 42102 705798
rect 41546 690618 42102 691174
rect 41546 654618 42102 655174
rect 41546 618618 42102 619174
rect 41546 582618 42102 583174
rect 41546 546618 42102 547174
rect 41546 510618 42102 511174
rect 41546 474618 42102 475174
rect 41546 438618 42102 439174
rect 41546 402618 42102 403174
rect 41546 366618 42102 367174
rect 41546 330618 42102 331174
rect 41546 294618 42102 295174
rect 41546 258618 42102 259174
rect 41546 222618 42102 223174
rect 41546 186618 42102 187174
rect 41546 150618 42102 151174
rect 41546 114618 42102 115174
rect 41546 78618 42102 79174
rect 41546 42618 42102 43174
rect 41546 6618 42102 7174
rect 41546 -1862 42102 -1306
rect 45266 706202 45822 706758
rect 45266 694338 45822 694894
rect 45266 658338 45822 658894
rect 45266 622338 45822 622894
rect 45266 586338 45822 586894
rect 45266 550338 45822 550894
rect 45266 514338 45822 514894
rect 45266 478338 45822 478894
rect 45266 442338 45822 442894
rect 45266 406338 45822 406894
rect 45266 370338 45822 370894
rect 45266 334338 45822 334894
rect 48986 707162 49542 707718
rect 48986 698058 49542 698614
rect 48986 662058 49542 662614
rect 48986 626058 49542 626614
rect 48986 590058 49542 590614
rect 48986 554058 49542 554614
rect 48986 518058 49542 518614
rect 48986 482058 49542 482614
rect 48986 446058 49542 446614
rect 48986 410058 49542 410614
rect 48986 374058 49542 374614
rect 48986 338058 49542 338614
rect 46970 327218 47206 327454
rect 46970 326898 47206 327134
rect 45266 298338 45822 298894
rect 48986 302058 49542 302614
rect 46970 291218 47206 291454
rect 46970 290898 47206 291134
rect 45266 262338 45822 262894
rect 48986 266058 49542 266614
rect 46970 255218 47206 255454
rect 46970 254898 47206 255134
rect 45266 226338 45822 226894
rect 48986 230058 49542 230614
rect 46970 219218 47206 219454
rect 46970 218898 47206 219134
rect 45266 190338 45822 190894
rect 48986 194058 49542 194614
rect 46970 183218 47206 183454
rect 46970 182898 47206 183134
rect 45266 154338 45822 154894
rect 48986 158058 49542 158614
rect 46970 147218 47206 147454
rect 46970 146898 47206 147134
rect 45266 118338 45822 118894
rect 48986 122058 49542 122614
rect 46970 111218 47206 111454
rect 46970 110898 47206 111134
rect 45266 82338 45822 82894
rect 48986 86058 49542 86614
rect 46970 75218 47206 75454
rect 46970 74898 47206 75134
rect 45266 46338 45822 46894
rect 48986 50058 49542 50614
rect 46970 39218 47206 39454
rect 46970 38898 47206 39134
rect 45266 10338 45822 10894
rect 45266 -2822 45822 -2266
rect 48986 14058 49542 14614
rect 48986 -3782 49542 -3226
rect 52706 708122 53262 708678
rect 52706 665778 53262 666334
rect 52706 629778 53262 630334
rect 52706 593778 53262 594334
rect 52706 557778 53262 558334
rect 52706 521778 53262 522334
rect 52706 485778 53262 486334
rect 52706 449778 53262 450334
rect 52706 413778 53262 414334
rect 52706 377778 53262 378334
rect 52706 341778 53262 342334
rect 52706 305778 53262 306334
rect 52706 269778 53262 270334
rect 52706 233778 53262 234334
rect 52706 197778 53262 198334
rect 52706 161778 53262 162334
rect 52706 125778 53262 126334
rect 52706 89778 53262 90334
rect 52706 53778 53262 54334
rect 52706 17778 53262 18334
rect 52706 -4742 53262 -4186
rect 56426 709082 56982 709638
rect 56426 669498 56982 670054
rect 56426 633498 56982 634054
rect 56426 597498 56982 598054
rect 56426 561498 56982 562054
rect 56426 525498 56982 526054
rect 56426 489498 56982 490054
rect 56426 453498 56982 454054
rect 56426 417498 56982 418054
rect 56426 381498 56982 382054
rect 56426 345498 56982 346054
rect 56426 309498 56982 310054
rect 56426 273498 56982 274054
rect 56426 237498 56982 238054
rect 56426 201498 56982 202054
rect 56426 165498 56982 166054
rect 56426 129498 56982 130054
rect 56426 93498 56982 94054
rect 56426 57498 56982 58054
rect 56426 21498 56982 22054
rect 56426 -5702 56982 -5146
rect 60146 710042 60702 710598
rect 60146 673218 60702 673774
rect 60146 637218 60702 637774
rect 60146 601218 60702 601774
rect 60146 565218 60702 565774
rect 60146 529218 60702 529774
rect 60146 493218 60702 493774
rect 60146 457218 60702 457774
rect 60146 421218 60702 421774
rect 60146 385218 60702 385774
rect 60146 349218 60702 349774
rect 63866 711002 64422 711558
rect 63866 676938 64422 677494
rect 63866 640938 64422 641494
rect 63866 604938 64422 605494
rect 63866 568938 64422 569494
rect 63866 532938 64422 533494
rect 63866 496938 64422 497494
rect 63866 460938 64422 461494
rect 63866 424938 64422 425494
rect 63866 388938 64422 389494
rect 63866 352938 64422 353494
rect 62330 330938 62566 331174
rect 62330 330618 62566 330854
rect 60146 313218 60702 313774
rect 63866 316938 64422 317494
rect 62330 294938 62566 295174
rect 62330 294618 62566 294854
rect 60146 277218 60702 277774
rect 63866 280938 64422 281494
rect 62330 258938 62566 259174
rect 62330 258618 62566 258854
rect 60146 241218 60702 241774
rect 63866 244938 64422 245494
rect 62330 222938 62566 223174
rect 62330 222618 62566 222854
rect 60146 205218 60702 205774
rect 63866 208938 64422 209494
rect 62330 186938 62566 187174
rect 62330 186618 62566 186854
rect 60146 169218 60702 169774
rect 63866 172938 64422 173494
rect 62330 150938 62566 151174
rect 62330 150618 62566 150854
rect 60146 133218 60702 133774
rect 63866 136938 64422 137494
rect 62330 114938 62566 115174
rect 62330 114618 62566 114854
rect 60146 97218 60702 97774
rect 63866 100938 64422 101494
rect 62330 78938 62566 79174
rect 62330 78618 62566 78854
rect 60146 61218 60702 61774
rect 63866 64938 64422 65494
rect 62330 42938 62566 43174
rect 62330 42618 62566 42854
rect 60146 25218 60702 25774
rect 63866 28938 64422 29494
rect 62330 6938 62566 7174
rect 62330 6618 62566 6854
rect 60146 -6662 60702 -6106
rect 63866 -7622 64422 -7066
rect 73826 704282 74382 704838
rect 73826 686898 74382 687454
rect 73826 650898 74382 651454
rect 73826 614898 74382 615454
rect 73826 578898 74382 579454
rect 73826 542898 74382 543454
rect 73826 506898 74382 507454
rect 73826 470898 74382 471454
rect 73826 434898 74382 435454
rect 73826 398898 74382 399454
rect 73826 362898 74382 363454
rect 77546 705242 78102 705798
rect 77546 690618 78102 691174
rect 77546 654618 78102 655174
rect 77546 618618 78102 619174
rect 77546 582618 78102 583174
rect 77546 546618 78102 547174
rect 77546 510618 78102 511174
rect 77546 474618 78102 475174
rect 77546 438618 78102 439174
rect 77546 402618 78102 403174
rect 77546 366618 78102 367174
rect 81266 706202 81822 706758
rect 81266 694338 81822 694894
rect 81266 658338 81822 658894
rect 81266 622338 81822 622894
rect 81266 586338 81822 586894
rect 81266 550338 81822 550894
rect 81266 514338 81822 514894
rect 81266 478338 81822 478894
rect 81266 442338 81822 442894
rect 81266 406338 81822 406894
rect 81266 370338 81822 370894
rect 81266 334338 81822 334894
rect 73826 326898 74382 327454
rect 77690 327218 77926 327454
rect 77690 326898 77926 327134
rect 81266 298338 81822 298894
rect 73826 290898 74382 291454
rect 77690 291218 77926 291454
rect 77690 290898 77926 291134
rect 81266 262338 81822 262894
rect 73826 254898 74382 255454
rect 77690 255218 77926 255454
rect 77690 254898 77926 255134
rect 81266 226338 81822 226894
rect 73826 218898 74382 219454
rect 77690 219218 77926 219454
rect 77690 218898 77926 219134
rect 81266 190338 81822 190894
rect 73826 182898 74382 183454
rect 77690 183218 77926 183454
rect 77690 182898 77926 183134
rect 81266 154338 81822 154894
rect 73826 146898 74382 147454
rect 77690 147218 77926 147454
rect 77690 146898 77926 147134
rect 81266 118338 81822 118894
rect 73826 110898 74382 111454
rect 77690 111218 77926 111454
rect 77690 110898 77926 111134
rect 81266 82338 81822 82894
rect 73826 74898 74382 75454
rect 77690 75218 77926 75454
rect 77690 74898 77926 75134
rect 81266 46338 81822 46894
rect 73826 38898 74382 39454
rect 77690 39218 77926 39454
rect 77690 38898 77926 39134
rect 73826 2898 74382 3454
rect 73826 -902 74382 -346
rect 81266 10338 81822 10894
rect 81266 -2822 81822 -2266
rect 84986 707162 85542 707718
rect 84986 698058 85542 698614
rect 84986 662058 85542 662614
rect 84986 626058 85542 626614
rect 84986 590058 85542 590614
rect 84986 554058 85542 554614
rect 84986 518058 85542 518614
rect 84986 482058 85542 482614
rect 84986 446058 85542 446614
rect 84986 410058 85542 410614
rect 84986 374058 85542 374614
rect 84986 338058 85542 338614
rect 84986 302058 85542 302614
rect 84986 266058 85542 266614
rect 84986 230058 85542 230614
rect 84986 194058 85542 194614
rect 84986 158058 85542 158614
rect 84986 122058 85542 122614
rect 84986 86058 85542 86614
rect 84986 50058 85542 50614
rect 84986 14058 85542 14614
rect 84986 -3782 85542 -3226
rect 88706 708122 89262 708678
rect 88706 665778 89262 666334
rect 88706 629778 89262 630334
rect 88706 593778 89262 594334
rect 88706 557778 89262 558334
rect 88706 521778 89262 522334
rect 88706 485778 89262 486334
rect 88706 449778 89262 450334
rect 88706 413778 89262 414334
rect 88706 377778 89262 378334
rect 92426 709082 92982 709638
rect 92426 669498 92982 670054
rect 92426 633498 92982 634054
rect 92426 597498 92982 598054
rect 92426 561498 92982 562054
rect 92426 525498 92982 526054
rect 92426 489498 92982 490054
rect 92426 453498 92982 454054
rect 92426 417498 92982 418054
rect 92426 381498 92982 382054
rect 96146 710042 96702 710598
rect 96146 673218 96702 673774
rect 96146 637218 96702 637774
rect 96146 601218 96702 601774
rect 96146 565218 96702 565774
rect 96146 529218 96702 529774
rect 96146 493218 96702 493774
rect 96146 457218 96702 457774
rect 96146 421218 96702 421774
rect 96146 385218 96702 385774
rect 88706 341778 89262 342334
rect 96146 349218 96702 349774
rect 93050 330938 93286 331174
rect 93050 330618 93286 330854
rect 88706 305778 89262 306334
rect 96146 313218 96702 313774
rect 93050 294938 93286 295174
rect 93050 294618 93286 294854
rect 88706 269778 89262 270334
rect 96146 277218 96702 277774
rect 93050 258938 93286 259174
rect 93050 258618 93286 258854
rect 88706 233778 89262 234334
rect 96146 241218 96702 241774
rect 93050 222938 93286 223174
rect 93050 222618 93286 222854
rect 88706 197778 89262 198334
rect 96146 205218 96702 205774
rect 93050 186938 93286 187174
rect 93050 186618 93286 186854
rect 88706 161778 89262 162334
rect 96146 169218 96702 169774
rect 93050 150938 93286 151174
rect 93050 150618 93286 150854
rect 88706 125778 89262 126334
rect 96146 133218 96702 133774
rect 93050 114938 93286 115174
rect 93050 114618 93286 114854
rect 88706 89778 89262 90334
rect 96146 97218 96702 97774
rect 93050 78938 93286 79174
rect 93050 78618 93286 78854
rect 88706 53778 89262 54334
rect 96146 61218 96702 61774
rect 93050 42938 93286 43174
rect 93050 42618 93286 42854
rect 88706 17778 89262 18334
rect 96146 25218 96702 25774
rect 93050 6938 93286 7174
rect 93050 6618 93286 6854
rect 88706 -4742 89262 -4186
rect 96146 -6662 96702 -6106
rect 99866 711002 100422 711558
rect 99866 676938 100422 677494
rect 99866 640938 100422 641494
rect 99866 604938 100422 605494
rect 99866 568938 100422 569494
rect 99866 532938 100422 533494
rect 99866 496938 100422 497494
rect 99866 460938 100422 461494
rect 99866 424938 100422 425494
rect 99866 388938 100422 389494
rect 99866 352938 100422 353494
rect 109826 704282 110382 704838
rect 109826 686898 110382 687454
rect 109826 650898 110382 651454
rect 109826 614898 110382 615454
rect 109826 578898 110382 579454
rect 109826 542898 110382 543454
rect 109826 506898 110382 507454
rect 109826 470898 110382 471454
rect 109826 434898 110382 435454
rect 109826 398898 110382 399454
rect 109826 362898 110382 363454
rect 108410 327218 108646 327454
rect 108410 326898 108646 327134
rect 109826 326898 110382 327454
rect 99866 316938 100422 317494
rect 108410 291218 108646 291454
rect 108410 290898 108646 291134
rect 109826 290898 110382 291454
rect 99866 280938 100422 281494
rect 108410 255218 108646 255454
rect 108410 254898 108646 255134
rect 109826 254898 110382 255454
rect 99866 244938 100422 245494
rect 108410 219218 108646 219454
rect 108410 218898 108646 219134
rect 109826 218898 110382 219454
rect 99866 208938 100422 209494
rect 108410 183218 108646 183454
rect 108410 182898 108646 183134
rect 109826 182898 110382 183454
rect 99866 172938 100422 173494
rect 108410 147218 108646 147454
rect 108410 146898 108646 147134
rect 109826 146898 110382 147454
rect 99866 136938 100422 137494
rect 108410 111218 108646 111454
rect 108410 110898 108646 111134
rect 109826 110898 110382 111454
rect 99866 100938 100422 101494
rect 108410 75218 108646 75454
rect 108410 74898 108646 75134
rect 109826 74898 110382 75454
rect 99866 64938 100422 65494
rect 108410 39218 108646 39454
rect 108410 38898 108646 39134
rect 109826 38898 110382 39454
rect 99866 28938 100422 29494
rect 99866 -7622 100422 -7066
rect 109826 2898 110382 3454
rect 109826 -902 110382 -346
rect 113546 705242 114102 705798
rect 113546 690618 114102 691174
rect 113546 654618 114102 655174
rect 113546 618618 114102 619174
rect 113546 582618 114102 583174
rect 113546 546618 114102 547174
rect 113546 510618 114102 511174
rect 113546 474618 114102 475174
rect 113546 438618 114102 439174
rect 113546 402618 114102 403174
rect 113546 366618 114102 367174
rect 113546 330618 114102 331174
rect 113546 294618 114102 295174
rect 113546 258618 114102 259174
rect 113546 222618 114102 223174
rect 113546 186618 114102 187174
rect 113546 150618 114102 151174
rect 113546 114618 114102 115174
rect 113546 78618 114102 79174
rect 113546 42618 114102 43174
rect 113546 6618 114102 7174
rect 113546 -1862 114102 -1306
rect 117266 706202 117822 706758
rect 117266 694338 117822 694894
rect 117266 658338 117822 658894
rect 117266 622338 117822 622894
rect 117266 586338 117822 586894
rect 117266 550338 117822 550894
rect 117266 514338 117822 514894
rect 117266 478338 117822 478894
rect 117266 442338 117822 442894
rect 117266 406338 117822 406894
rect 117266 370338 117822 370894
rect 117266 334338 117822 334894
rect 117266 298338 117822 298894
rect 117266 262338 117822 262894
rect 117266 226338 117822 226894
rect 117266 190338 117822 190894
rect 117266 154338 117822 154894
rect 117266 118338 117822 118894
rect 117266 82338 117822 82894
rect 117266 46338 117822 46894
rect 117266 10338 117822 10894
rect 117266 -2822 117822 -2266
rect 120986 707162 121542 707718
rect 120986 698058 121542 698614
rect 120986 662058 121542 662614
rect 120986 626058 121542 626614
rect 120986 590058 121542 590614
rect 120986 554058 121542 554614
rect 120986 518058 121542 518614
rect 120986 482058 121542 482614
rect 120986 446058 121542 446614
rect 120986 410058 121542 410614
rect 120986 374058 121542 374614
rect 120986 338058 121542 338614
rect 124706 708122 125262 708678
rect 124706 665778 125262 666334
rect 124706 629778 125262 630334
rect 124706 593778 125262 594334
rect 124706 557778 125262 558334
rect 124706 521778 125262 522334
rect 124706 485778 125262 486334
rect 124706 449778 125262 450334
rect 124706 413778 125262 414334
rect 124706 377778 125262 378334
rect 124706 341778 125262 342334
rect 123770 330938 124006 331174
rect 123770 330618 124006 330854
rect 120986 302058 121542 302614
rect 124706 305778 125262 306334
rect 123770 294938 124006 295174
rect 123770 294618 124006 294854
rect 120986 266058 121542 266614
rect 124706 269778 125262 270334
rect 123770 258938 124006 259174
rect 123770 258618 124006 258854
rect 120986 230058 121542 230614
rect 124706 233778 125262 234334
rect 123770 222938 124006 223174
rect 123770 222618 124006 222854
rect 120986 194058 121542 194614
rect 124706 197778 125262 198334
rect 123770 186938 124006 187174
rect 123770 186618 124006 186854
rect 120986 158058 121542 158614
rect 124706 161778 125262 162334
rect 123770 150938 124006 151174
rect 123770 150618 124006 150854
rect 120986 122058 121542 122614
rect 124706 125778 125262 126334
rect 123770 114938 124006 115174
rect 123770 114618 124006 114854
rect 120986 86058 121542 86614
rect 124706 89778 125262 90334
rect 123770 78938 124006 79174
rect 123770 78618 124006 78854
rect 120986 50058 121542 50614
rect 124706 53778 125262 54334
rect 123770 42938 124006 43174
rect 123770 42618 124006 42854
rect 120986 14058 121542 14614
rect 124706 17778 125262 18334
rect 123770 6938 124006 7174
rect 123770 6618 124006 6854
rect 120986 -3782 121542 -3226
rect 124706 -4742 125262 -4186
rect 128426 709082 128982 709638
rect 128426 669498 128982 670054
rect 128426 633498 128982 634054
rect 128426 597498 128982 598054
rect 128426 561498 128982 562054
rect 128426 525498 128982 526054
rect 128426 489498 128982 490054
rect 128426 453498 128982 454054
rect 128426 417498 128982 418054
rect 128426 381498 128982 382054
rect 128426 345498 128982 346054
rect 128426 309498 128982 310054
rect 128426 273498 128982 274054
rect 128426 237498 128982 238054
rect 128426 201498 128982 202054
rect 128426 165498 128982 166054
rect 128426 129498 128982 130054
rect 128426 93498 128982 94054
rect 128426 57498 128982 58054
rect 128426 21498 128982 22054
rect 128426 -5702 128982 -5146
rect 132146 710042 132702 710598
rect 132146 673218 132702 673774
rect 132146 637218 132702 637774
rect 132146 601218 132702 601774
rect 132146 565218 132702 565774
rect 132146 529218 132702 529774
rect 132146 493218 132702 493774
rect 132146 457218 132702 457774
rect 132146 421218 132702 421774
rect 132146 385218 132702 385774
rect 132146 349218 132702 349774
rect 132146 313218 132702 313774
rect 132146 277218 132702 277774
rect 132146 241218 132702 241774
rect 132146 205218 132702 205774
rect 132146 169218 132702 169774
rect 132146 133218 132702 133774
rect 132146 97218 132702 97774
rect 132146 61218 132702 61774
rect 132146 25218 132702 25774
rect 132146 -6662 132702 -6106
rect 135866 711002 136422 711558
rect 135866 676938 136422 677494
rect 135866 640938 136422 641494
rect 135866 604938 136422 605494
rect 135866 568938 136422 569494
rect 135866 532938 136422 533494
rect 135866 496938 136422 497494
rect 135866 460938 136422 461494
rect 135866 424938 136422 425494
rect 135866 388938 136422 389494
rect 135866 352938 136422 353494
rect 145826 704282 146382 704838
rect 145826 686898 146382 687454
rect 145826 650898 146382 651454
rect 145826 614898 146382 615454
rect 145826 578898 146382 579454
rect 145826 542898 146382 543454
rect 145826 506898 146382 507454
rect 145826 470898 146382 471454
rect 145826 434898 146382 435454
rect 145826 398898 146382 399454
rect 145826 362898 146382 363454
rect 139130 327218 139366 327454
rect 139130 326898 139366 327134
rect 145826 326898 146382 327454
rect 135866 316938 136422 317494
rect 139130 291218 139366 291454
rect 139130 290898 139366 291134
rect 145826 290898 146382 291454
rect 135866 280938 136422 281494
rect 139130 255218 139366 255454
rect 139130 254898 139366 255134
rect 145826 254898 146382 255454
rect 135866 244938 136422 245494
rect 139130 219218 139366 219454
rect 139130 218898 139366 219134
rect 145826 218898 146382 219454
rect 135866 208938 136422 209494
rect 139130 183218 139366 183454
rect 139130 182898 139366 183134
rect 145826 182898 146382 183454
rect 135866 172938 136422 173494
rect 139130 147218 139366 147454
rect 139130 146898 139366 147134
rect 145826 146898 146382 147454
rect 135866 136938 136422 137494
rect 139130 111218 139366 111454
rect 139130 110898 139366 111134
rect 145826 110898 146382 111454
rect 135866 100938 136422 101494
rect 139130 75218 139366 75454
rect 139130 74898 139366 75134
rect 145826 74898 146382 75454
rect 135866 64938 136422 65494
rect 139130 39218 139366 39454
rect 139130 38898 139366 39134
rect 145826 38898 146382 39454
rect 135866 28938 136422 29494
rect 135866 -7622 136422 -7066
rect 145826 2898 146382 3454
rect 145826 -902 146382 -346
rect 149546 705242 150102 705798
rect 149546 690618 150102 691174
rect 149546 654618 150102 655174
rect 149546 618618 150102 619174
rect 149546 582618 150102 583174
rect 149546 546618 150102 547174
rect 149546 510618 150102 511174
rect 149546 474618 150102 475174
rect 149546 438618 150102 439174
rect 149546 402618 150102 403174
rect 149546 366618 150102 367174
rect 149546 330618 150102 331174
rect 149546 294618 150102 295174
rect 149546 258618 150102 259174
rect 149546 222618 150102 223174
rect 149546 186618 150102 187174
rect 149546 150618 150102 151174
rect 149546 114618 150102 115174
rect 149546 78618 150102 79174
rect 149546 42618 150102 43174
rect 149546 6618 150102 7174
rect 149546 -1862 150102 -1306
rect 153266 706202 153822 706758
rect 153266 694338 153822 694894
rect 153266 658338 153822 658894
rect 153266 622338 153822 622894
rect 153266 586338 153822 586894
rect 153266 550338 153822 550894
rect 153266 514338 153822 514894
rect 153266 478338 153822 478894
rect 153266 442338 153822 442894
rect 153266 406338 153822 406894
rect 153266 370338 153822 370894
rect 153266 334338 153822 334894
rect 156986 707162 157542 707718
rect 156986 698058 157542 698614
rect 156986 662058 157542 662614
rect 156986 626058 157542 626614
rect 156986 590058 157542 590614
rect 156986 554058 157542 554614
rect 156986 518058 157542 518614
rect 156986 482058 157542 482614
rect 156986 446058 157542 446614
rect 156986 410058 157542 410614
rect 156986 374058 157542 374614
rect 156986 338058 157542 338614
rect 154490 330938 154726 331174
rect 154490 330618 154726 330854
rect 153266 298338 153822 298894
rect 156986 302058 157542 302614
rect 154490 294938 154726 295174
rect 154490 294618 154726 294854
rect 153266 262338 153822 262894
rect 156986 266058 157542 266614
rect 154490 258938 154726 259174
rect 154490 258618 154726 258854
rect 153266 226338 153822 226894
rect 156986 230058 157542 230614
rect 154490 222938 154726 223174
rect 154490 222618 154726 222854
rect 153266 190338 153822 190894
rect 156986 194058 157542 194614
rect 154490 186938 154726 187174
rect 154490 186618 154726 186854
rect 153266 154338 153822 154894
rect 156986 158058 157542 158614
rect 154490 150938 154726 151174
rect 154490 150618 154726 150854
rect 153266 118338 153822 118894
rect 156986 122058 157542 122614
rect 154490 114938 154726 115174
rect 154490 114618 154726 114854
rect 153266 82338 153822 82894
rect 156986 86058 157542 86614
rect 154490 78938 154726 79174
rect 154490 78618 154726 78854
rect 153266 46338 153822 46894
rect 156986 50058 157542 50614
rect 154490 42938 154726 43174
rect 154490 42618 154726 42854
rect 153266 10338 153822 10894
rect 156986 14058 157542 14614
rect 154490 6938 154726 7174
rect 154490 6618 154726 6854
rect 153266 -2822 153822 -2266
rect 156986 -3782 157542 -3226
rect 160706 708122 161262 708678
rect 160706 665778 161262 666334
rect 160706 629778 161262 630334
rect 160706 593778 161262 594334
rect 160706 557778 161262 558334
rect 160706 521778 161262 522334
rect 160706 485778 161262 486334
rect 160706 449778 161262 450334
rect 160706 413778 161262 414334
rect 160706 377778 161262 378334
rect 160706 341778 161262 342334
rect 160706 305778 161262 306334
rect 160706 269778 161262 270334
rect 160706 233778 161262 234334
rect 160706 197778 161262 198334
rect 160706 161778 161262 162334
rect 160706 125778 161262 126334
rect 160706 89778 161262 90334
rect 160706 53778 161262 54334
rect 160706 17778 161262 18334
rect 160706 -4742 161262 -4186
rect 164426 709082 164982 709638
rect 164426 669498 164982 670054
rect 164426 633498 164982 634054
rect 164426 597498 164982 598054
rect 164426 561498 164982 562054
rect 164426 525498 164982 526054
rect 164426 489498 164982 490054
rect 164426 453498 164982 454054
rect 164426 417498 164982 418054
rect 164426 381498 164982 382054
rect 164426 345498 164982 346054
rect 164426 309498 164982 310054
rect 164426 273498 164982 274054
rect 164426 237498 164982 238054
rect 164426 201498 164982 202054
rect 164426 165498 164982 166054
rect 164426 129498 164982 130054
rect 164426 93498 164982 94054
rect 164426 57498 164982 58054
rect 164426 21498 164982 22054
rect 164426 -5702 164982 -5146
rect 168146 710042 168702 710598
rect 168146 673218 168702 673774
rect 168146 637218 168702 637774
rect 168146 601218 168702 601774
rect 168146 565218 168702 565774
rect 168146 529218 168702 529774
rect 168146 493218 168702 493774
rect 168146 457218 168702 457774
rect 168146 421218 168702 421774
rect 168146 385218 168702 385774
rect 168146 349218 168702 349774
rect 171866 711002 172422 711558
rect 171866 676938 172422 677494
rect 171866 640938 172422 641494
rect 171866 604938 172422 605494
rect 171866 568938 172422 569494
rect 171866 532938 172422 533494
rect 171866 496938 172422 497494
rect 171866 460938 172422 461494
rect 171866 424938 172422 425494
rect 171866 388938 172422 389494
rect 171866 352938 172422 353494
rect 169850 327218 170086 327454
rect 169850 326898 170086 327134
rect 168146 313218 168702 313774
rect 171866 316938 172422 317494
rect 169850 291218 170086 291454
rect 169850 290898 170086 291134
rect 168146 277218 168702 277774
rect 171866 280938 172422 281494
rect 169850 255218 170086 255454
rect 169850 254898 170086 255134
rect 168146 241218 168702 241774
rect 171866 244938 172422 245494
rect 169850 219218 170086 219454
rect 169850 218898 170086 219134
rect 168146 205218 168702 205774
rect 171866 208938 172422 209494
rect 169850 183218 170086 183454
rect 169850 182898 170086 183134
rect 168146 169218 168702 169774
rect 171866 172938 172422 173494
rect 169850 147218 170086 147454
rect 169850 146898 170086 147134
rect 168146 133218 168702 133774
rect 171866 136938 172422 137494
rect 169850 111218 170086 111454
rect 169850 110898 170086 111134
rect 168146 97218 168702 97774
rect 171866 100938 172422 101494
rect 169850 75218 170086 75454
rect 169850 74898 170086 75134
rect 168146 61218 168702 61774
rect 171866 64938 172422 65494
rect 169850 39218 170086 39454
rect 169850 38898 170086 39134
rect 168146 25218 168702 25774
rect 168146 -6662 168702 -6106
rect 171866 28938 172422 29494
rect 171866 -7622 172422 -7066
rect 181826 704282 182382 704838
rect 181826 686898 182382 687454
rect 181826 650898 182382 651454
rect 181826 614898 182382 615454
rect 181826 578898 182382 579454
rect 181826 542898 182382 543454
rect 181826 506898 182382 507454
rect 181826 470898 182382 471454
rect 181826 434898 182382 435454
rect 181826 398898 182382 399454
rect 181826 362898 182382 363454
rect 185546 705242 186102 705798
rect 185546 690618 186102 691174
rect 185546 654618 186102 655174
rect 185546 618618 186102 619174
rect 185546 582618 186102 583174
rect 185546 546618 186102 547174
rect 185546 510618 186102 511174
rect 185546 474618 186102 475174
rect 185546 438618 186102 439174
rect 185546 402618 186102 403174
rect 185546 366618 186102 367174
rect 189266 706202 189822 706758
rect 189266 694338 189822 694894
rect 189266 658338 189822 658894
rect 189266 622338 189822 622894
rect 189266 586338 189822 586894
rect 189266 550338 189822 550894
rect 189266 514338 189822 514894
rect 189266 478338 189822 478894
rect 189266 442338 189822 442894
rect 189266 406338 189822 406894
rect 189266 370338 189822 370894
rect 189266 334338 189822 334894
rect 185210 330938 185446 331174
rect 185210 330618 185446 330854
rect 181826 326898 182382 327454
rect 189266 298338 189822 298894
rect 185210 294938 185446 295174
rect 185210 294618 185446 294854
rect 181826 290898 182382 291454
rect 189266 262338 189822 262894
rect 185210 258938 185446 259174
rect 185210 258618 185446 258854
rect 181826 254898 182382 255454
rect 189266 226338 189822 226894
rect 185210 222938 185446 223174
rect 185210 222618 185446 222854
rect 181826 218898 182382 219454
rect 189266 190338 189822 190894
rect 185210 186938 185446 187174
rect 185210 186618 185446 186854
rect 181826 182898 182382 183454
rect 189266 154338 189822 154894
rect 185210 150938 185446 151174
rect 185210 150618 185446 150854
rect 181826 146898 182382 147454
rect 189266 118338 189822 118894
rect 185210 114938 185446 115174
rect 185210 114618 185446 114854
rect 181826 110898 182382 111454
rect 189266 82338 189822 82894
rect 185210 78938 185446 79174
rect 185210 78618 185446 78854
rect 181826 74898 182382 75454
rect 189266 46338 189822 46894
rect 185210 42938 185446 43174
rect 185210 42618 185446 42854
rect 181826 38898 182382 39454
rect 189266 10338 189822 10894
rect 185210 6938 185446 7174
rect 185210 6618 185446 6854
rect 181826 2898 182382 3454
rect 181826 -902 182382 -346
rect 189266 -2822 189822 -2266
rect 192986 707162 193542 707718
rect 192986 698058 193542 698614
rect 192986 662058 193542 662614
rect 192986 626058 193542 626614
rect 192986 590058 193542 590614
rect 192986 554058 193542 554614
rect 192986 518058 193542 518614
rect 192986 482058 193542 482614
rect 192986 446058 193542 446614
rect 192986 410058 193542 410614
rect 192986 374058 193542 374614
rect 192986 338058 193542 338614
rect 192986 302058 193542 302614
rect 192986 266058 193542 266614
rect 192986 230058 193542 230614
rect 192986 194058 193542 194614
rect 192986 158058 193542 158614
rect 192986 122058 193542 122614
rect 192986 86058 193542 86614
rect 192986 50058 193542 50614
rect 192986 14058 193542 14614
rect 192986 -3782 193542 -3226
rect 196706 708122 197262 708678
rect 196706 665778 197262 666334
rect 196706 629778 197262 630334
rect 196706 593778 197262 594334
rect 196706 557778 197262 558334
rect 196706 521778 197262 522334
rect 196706 485778 197262 486334
rect 196706 449778 197262 450334
rect 196706 413778 197262 414334
rect 196706 377778 197262 378334
rect 200426 709082 200982 709638
rect 200426 669498 200982 670054
rect 200426 633498 200982 634054
rect 200426 597498 200982 598054
rect 200426 561498 200982 562054
rect 200426 525498 200982 526054
rect 200426 489498 200982 490054
rect 200426 453498 200982 454054
rect 200426 417498 200982 418054
rect 200426 381498 200982 382054
rect 204146 710042 204702 710598
rect 204146 673218 204702 673774
rect 204146 637218 204702 637774
rect 204146 601218 204702 601774
rect 204146 565218 204702 565774
rect 204146 529218 204702 529774
rect 204146 493218 204702 493774
rect 204146 457218 204702 457774
rect 204146 421218 204702 421774
rect 204146 385218 204702 385774
rect 196706 341778 197262 342334
rect 204146 349218 204702 349774
rect 200570 327218 200806 327454
rect 200570 326898 200806 327134
rect 196706 305778 197262 306334
rect 204146 313218 204702 313774
rect 200570 291218 200806 291454
rect 200570 290898 200806 291134
rect 196706 269778 197262 270334
rect 204146 277218 204702 277774
rect 200570 255218 200806 255454
rect 200570 254898 200806 255134
rect 196706 233778 197262 234334
rect 204146 241218 204702 241774
rect 200570 219218 200806 219454
rect 200570 218898 200806 219134
rect 196706 197778 197262 198334
rect 204146 205218 204702 205774
rect 200570 183218 200806 183454
rect 200570 182898 200806 183134
rect 196706 161778 197262 162334
rect 204146 169218 204702 169774
rect 200570 147218 200806 147454
rect 200570 146898 200806 147134
rect 196706 125778 197262 126334
rect 204146 133218 204702 133774
rect 200570 111218 200806 111454
rect 200570 110898 200806 111134
rect 196706 89778 197262 90334
rect 204146 97218 204702 97774
rect 200570 75218 200806 75454
rect 200570 74898 200806 75134
rect 196706 53778 197262 54334
rect 204146 61218 204702 61774
rect 200570 39218 200806 39454
rect 200570 38898 200806 39134
rect 196706 17778 197262 18334
rect 196706 -4742 197262 -4186
rect 204146 25218 204702 25774
rect 204146 -6662 204702 -6106
rect 207866 711002 208422 711558
rect 207866 676938 208422 677494
rect 207866 640938 208422 641494
rect 207866 604938 208422 605494
rect 207866 568938 208422 569494
rect 207866 532938 208422 533494
rect 207866 496938 208422 497494
rect 207866 460938 208422 461494
rect 207866 424938 208422 425494
rect 207866 388938 208422 389494
rect 207866 352938 208422 353494
rect 217826 704282 218382 704838
rect 217826 686898 218382 687454
rect 217826 650898 218382 651454
rect 217826 614898 218382 615454
rect 217826 578898 218382 579454
rect 217826 542898 218382 543454
rect 217826 506898 218382 507454
rect 217826 470898 218382 471454
rect 217826 434898 218382 435454
rect 217826 398898 218382 399454
rect 217826 362898 218382 363454
rect 215930 330938 216166 331174
rect 215930 330618 216166 330854
rect 207866 316938 208422 317494
rect 217826 326898 218382 327454
rect 215930 294938 216166 295174
rect 215930 294618 216166 294854
rect 207866 280938 208422 281494
rect 217826 290898 218382 291454
rect 215930 258938 216166 259174
rect 215930 258618 216166 258854
rect 207866 244938 208422 245494
rect 217826 254898 218382 255454
rect 215930 222938 216166 223174
rect 215930 222618 216166 222854
rect 207866 208938 208422 209494
rect 217826 218898 218382 219454
rect 215930 186938 216166 187174
rect 215930 186618 216166 186854
rect 207866 172938 208422 173494
rect 217826 182898 218382 183454
rect 215930 150938 216166 151174
rect 215930 150618 216166 150854
rect 207866 136938 208422 137494
rect 217826 146898 218382 147454
rect 215930 114938 216166 115174
rect 215930 114618 216166 114854
rect 207866 100938 208422 101494
rect 217826 110898 218382 111454
rect 215930 78938 216166 79174
rect 215930 78618 216166 78854
rect 207866 64938 208422 65494
rect 217826 74898 218382 75454
rect 215930 42938 216166 43174
rect 215930 42618 216166 42854
rect 207866 28938 208422 29494
rect 217826 38898 218382 39454
rect 215930 6938 216166 7174
rect 215930 6618 216166 6854
rect 207866 -7622 208422 -7066
rect 217826 2898 218382 3454
rect 217826 -902 218382 -346
rect 221546 705242 222102 705798
rect 221546 690618 222102 691174
rect 221546 654618 222102 655174
rect 221546 618618 222102 619174
rect 221546 582618 222102 583174
rect 221546 546618 222102 547174
rect 221546 510618 222102 511174
rect 221546 474618 222102 475174
rect 221546 438618 222102 439174
rect 221546 402618 222102 403174
rect 221546 366618 222102 367174
rect 221546 330618 222102 331174
rect 221546 294618 222102 295174
rect 221546 258618 222102 259174
rect 221546 222618 222102 223174
rect 221546 186618 222102 187174
rect 221546 150618 222102 151174
rect 221546 114618 222102 115174
rect 221546 78618 222102 79174
rect 221546 42618 222102 43174
rect 221546 6618 222102 7174
rect 221546 -1862 222102 -1306
rect 225266 706202 225822 706758
rect 225266 694338 225822 694894
rect 225266 658338 225822 658894
rect 225266 622338 225822 622894
rect 225266 586338 225822 586894
rect 225266 550338 225822 550894
rect 225266 514338 225822 514894
rect 225266 478338 225822 478894
rect 225266 442338 225822 442894
rect 225266 406338 225822 406894
rect 225266 370338 225822 370894
rect 225266 334338 225822 334894
rect 225266 298338 225822 298894
rect 225266 262338 225822 262894
rect 225266 226338 225822 226894
rect 225266 190338 225822 190894
rect 225266 154338 225822 154894
rect 225266 118338 225822 118894
rect 225266 82338 225822 82894
rect 225266 46338 225822 46894
rect 225266 10338 225822 10894
rect 225266 -2822 225822 -2266
rect 228986 707162 229542 707718
rect 228986 698058 229542 698614
rect 228986 662058 229542 662614
rect 228986 626058 229542 626614
rect 228986 590058 229542 590614
rect 228986 554058 229542 554614
rect 228986 518058 229542 518614
rect 228986 482058 229542 482614
rect 228986 446058 229542 446614
rect 228986 410058 229542 410614
rect 228986 374058 229542 374614
rect 228986 338058 229542 338614
rect 232706 708122 233262 708678
rect 232706 665778 233262 666334
rect 232706 629778 233262 630334
rect 232706 593778 233262 594334
rect 232706 557778 233262 558334
rect 232706 521778 233262 522334
rect 232706 485778 233262 486334
rect 232706 449778 233262 450334
rect 232706 413778 233262 414334
rect 232706 377778 233262 378334
rect 232706 341778 233262 342334
rect 231290 327218 231526 327454
rect 231290 326898 231526 327134
rect 228986 302058 229542 302614
rect 232706 305778 233262 306334
rect 231290 291218 231526 291454
rect 231290 290898 231526 291134
rect 228986 266058 229542 266614
rect 232706 269778 233262 270334
rect 231290 255218 231526 255454
rect 231290 254898 231526 255134
rect 228986 230058 229542 230614
rect 232706 233778 233262 234334
rect 231290 219218 231526 219454
rect 231290 218898 231526 219134
rect 228986 194058 229542 194614
rect 232706 197778 233262 198334
rect 231290 183218 231526 183454
rect 231290 182898 231526 183134
rect 228986 158058 229542 158614
rect 232706 161778 233262 162334
rect 231290 147218 231526 147454
rect 231290 146898 231526 147134
rect 228986 122058 229542 122614
rect 232706 125778 233262 126334
rect 231290 111218 231526 111454
rect 231290 110898 231526 111134
rect 228986 86058 229542 86614
rect 232706 89778 233262 90334
rect 231290 75218 231526 75454
rect 231290 74898 231526 75134
rect 228986 50058 229542 50614
rect 232706 53778 233262 54334
rect 231290 39218 231526 39454
rect 231290 38898 231526 39134
rect 228986 14058 229542 14614
rect 228986 -3782 229542 -3226
rect 232706 17778 233262 18334
rect 232706 -4742 233262 -4186
rect 236426 709082 236982 709638
rect 236426 669498 236982 670054
rect 236426 633498 236982 634054
rect 236426 597498 236982 598054
rect 236426 561498 236982 562054
rect 236426 525498 236982 526054
rect 236426 489498 236982 490054
rect 236426 453498 236982 454054
rect 236426 417498 236982 418054
rect 236426 381498 236982 382054
rect 236426 345498 236982 346054
rect 236426 309498 236982 310054
rect 236426 273498 236982 274054
rect 236426 237498 236982 238054
rect 236426 201498 236982 202054
rect 236426 165498 236982 166054
rect 236426 129498 236982 130054
rect 236426 93498 236982 94054
rect 236426 57498 236982 58054
rect 240146 710042 240702 710598
rect 240146 673218 240702 673774
rect 240146 637218 240702 637774
rect 240146 601218 240702 601774
rect 240146 565218 240702 565774
rect 240146 529218 240702 529774
rect 240146 493218 240702 493774
rect 240146 457218 240702 457774
rect 240146 421218 240702 421774
rect 240146 385218 240702 385774
rect 240146 349218 240702 349774
rect 240146 313218 240702 313774
rect 240146 277218 240702 277774
rect 240146 241218 240702 241774
rect 240146 205218 240702 205774
rect 240146 169218 240702 169774
rect 240146 133218 240702 133774
rect 240146 97218 240702 97774
rect 240146 61218 240702 61774
rect 243866 711002 244422 711558
rect 243866 676938 244422 677494
rect 243866 640938 244422 641494
rect 243866 604938 244422 605494
rect 243866 568938 244422 569494
rect 243866 532938 244422 533494
rect 243866 496938 244422 497494
rect 243866 460938 244422 461494
rect 243866 424938 244422 425494
rect 243866 388938 244422 389494
rect 243866 352938 244422 353494
rect 253826 704282 254382 704838
rect 253826 686898 254382 687454
rect 253826 650898 254382 651454
rect 253826 614898 254382 615454
rect 253826 578898 254382 579454
rect 253826 542898 254382 543454
rect 253826 506898 254382 507454
rect 253826 470898 254382 471454
rect 253826 434898 254382 435454
rect 253826 398898 254382 399454
rect 253826 362898 254382 363454
rect 246650 330938 246886 331174
rect 246650 330618 246886 330854
rect 243866 316938 244422 317494
rect 253826 326898 254382 327454
rect 246650 294938 246886 295174
rect 246650 294618 246886 294854
rect 243866 280938 244422 281494
rect 253826 290898 254382 291454
rect 246650 258938 246886 259174
rect 246650 258618 246886 258854
rect 243866 244938 244422 245494
rect 253826 254898 254382 255454
rect 246650 222938 246886 223174
rect 246650 222618 246886 222854
rect 243866 208938 244422 209494
rect 253826 218898 254382 219454
rect 246650 186938 246886 187174
rect 246650 186618 246886 186854
rect 243866 172938 244422 173494
rect 253826 182898 254382 183454
rect 246650 150938 246886 151174
rect 246650 150618 246886 150854
rect 243866 136938 244422 137494
rect 253826 146898 254382 147454
rect 246650 114938 246886 115174
rect 246650 114618 246886 114854
rect 243866 100938 244422 101494
rect 253826 110898 254382 111454
rect 246650 78938 246886 79174
rect 246650 78618 246886 78854
rect 243866 64938 244422 65494
rect 253826 74898 254382 75454
rect 246650 42938 246886 43174
rect 246650 42618 246886 42854
rect 243866 28938 244422 29494
rect 253826 38898 254382 39454
rect 257546 705242 258102 705798
rect 257546 690618 258102 691174
rect 257546 654618 258102 655174
rect 257546 618618 258102 619174
rect 257546 582618 258102 583174
rect 257546 546618 258102 547174
rect 257546 510618 258102 511174
rect 257546 474618 258102 475174
rect 257546 438618 258102 439174
rect 257546 402618 258102 403174
rect 257546 366618 258102 367174
rect 257546 330618 258102 331174
rect 257546 294618 258102 295174
rect 257546 258618 258102 259174
rect 257546 222618 258102 223174
rect 257546 186618 258102 187174
rect 257546 150618 258102 151174
rect 257546 114618 258102 115174
rect 257546 78618 258102 79174
rect 257546 42618 258102 43174
rect 261266 706202 261822 706758
rect 261266 694338 261822 694894
rect 261266 658338 261822 658894
rect 261266 622338 261822 622894
rect 261266 586338 261822 586894
rect 261266 550338 261822 550894
rect 261266 514338 261822 514894
rect 261266 478338 261822 478894
rect 261266 442338 261822 442894
rect 261266 406338 261822 406894
rect 261266 370338 261822 370894
rect 261266 334338 261822 334894
rect 264986 707162 265542 707718
rect 264986 698058 265542 698614
rect 264986 662058 265542 662614
rect 264986 626058 265542 626614
rect 264986 590058 265542 590614
rect 264986 554058 265542 554614
rect 264986 518058 265542 518614
rect 264986 482058 265542 482614
rect 264986 446058 265542 446614
rect 264986 410058 265542 410614
rect 264986 374058 265542 374614
rect 264986 338058 265542 338614
rect 262010 327218 262246 327454
rect 262010 326898 262246 327134
rect 261266 298338 261822 298894
rect 264986 302058 265542 302614
rect 262010 291218 262246 291454
rect 262010 290898 262246 291134
rect 261266 262338 261822 262894
rect 264986 266058 265542 266614
rect 262010 255218 262246 255454
rect 262010 254898 262246 255134
rect 261266 226338 261822 226894
rect 264986 230058 265542 230614
rect 262010 219218 262246 219454
rect 262010 218898 262246 219134
rect 261266 190338 261822 190894
rect 264986 194058 265542 194614
rect 262010 183218 262246 183454
rect 262010 182898 262246 183134
rect 261266 154338 261822 154894
rect 264986 158058 265542 158614
rect 262010 147218 262246 147454
rect 262010 146898 262246 147134
rect 261266 118338 261822 118894
rect 264986 122058 265542 122614
rect 262010 111218 262246 111454
rect 262010 110898 262246 111134
rect 261266 82338 261822 82894
rect 264986 86058 265542 86614
rect 262010 75218 262246 75454
rect 262010 74898 262246 75134
rect 261266 46338 261822 46894
rect 236426 21498 236982 22054
rect 264986 50058 265542 50614
rect 262010 39218 262246 39454
rect 262010 38898 262246 39134
rect 261266 10338 261822 10894
rect 246650 6938 246886 7174
rect 246650 6618 246886 6854
rect 236426 -5702 236982 -5146
rect 253826 2898 254382 3454
rect 253826 -902 254382 -346
rect 261266 -2822 261822 -2266
rect 264986 14058 265542 14614
rect 264986 -3782 265542 -3226
rect 268706 708122 269262 708678
rect 268706 665778 269262 666334
rect 268706 629778 269262 630334
rect 268706 593778 269262 594334
rect 268706 557778 269262 558334
rect 268706 521778 269262 522334
rect 268706 485778 269262 486334
rect 268706 449778 269262 450334
rect 268706 413778 269262 414334
rect 268706 377778 269262 378334
rect 268706 341778 269262 342334
rect 268706 305778 269262 306334
rect 268706 269778 269262 270334
rect 268706 233778 269262 234334
rect 268706 197778 269262 198334
rect 268706 161778 269262 162334
rect 268706 125778 269262 126334
rect 268706 89778 269262 90334
rect 268706 53778 269262 54334
rect 268706 17778 269262 18334
rect 268706 -4742 269262 -4186
rect 272426 709082 272982 709638
rect 272426 669498 272982 670054
rect 272426 633498 272982 634054
rect 272426 597498 272982 598054
rect 272426 561498 272982 562054
rect 272426 525498 272982 526054
rect 272426 489498 272982 490054
rect 272426 453498 272982 454054
rect 272426 417498 272982 418054
rect 272426 381498 272982 382054
rect 272426 345498 272982 346054
rect 272426 309498 272982 310054
rect 272426 273498 272982 274054
rect 272426 237498 272982 238054
rect 272426 201498 272982 202054
rect 272426 165498 272982 166054
rect 272426 129498 272982 130054
rect 272426 93498 272982 94054
rect 272426 57498 272982 58054
rect 272426 21498 272982 22054
rect 272426 -5702 272982 -5146
rect 276146 710042 276702 710598
rect 276146 673218 276702 673774
rect 276146 637218 276702 637774
rect 276146 601218 276702 601774
rect 276146 565218 276702 565774
rect 276146 529218 276702 529774
rect 276146 493218 276702 493774
rect 276146 457218 276702 457774
rect 276146 421218 276702 421774
rect 276146 385218 276702 385774
rect 276146 349218 276702 349774
rect 279866 711002 280422 711558
rect 279866 676938 280422 677494
rect 279866 640938 280422 641494
rect 279866 604938 280422 605494
rect 279866 568938 280422 569494
rect 279866 532938 280422 533494
rect 279866 496938 280422 497494
rect 279866 460938 280422 461494
rect 279866 424938 280422 425494
rect 279866 388938 280422 389494
rect 279866 352938 280422 353494
rect 277370 330938 277606 331174
rect 277370 330618 277606 330854
rect 276146 313218 276702 313774
rect 279866 316938 280422 317494
rect 277370 294938 277606 295174
rect 277370 294618 277606 294854
rect 276146 277218 276702 277774
rect 279866 280938 280422 281494
rect 277370 258938 277606 259174
rect 277370 258618 277606 258854
rect 276146 241218 276702 241774
rect 279866 244938 280422 245494
rect 277370 222938 277606 223174
rect 277370 222618 277606 222854
rect 276146 205218 276702 205774
rect 279866 208938 280422 209494
rect 277370 186938 277606 187174
rect 277370 186618 277606 186854
rect 276146 169218 276702 169774
rect 279866 172938 280422 173494
rect 277370 150938 277606 151174
rect 277370 150618 277606 150854
rect 276146 133218 276702 133774
rect 279866 136938 280422 137494
rect 277370 114938 277606 115174
rect 277370 114618 277606 114854
rect 276146 97218 276702 97774
rect 279866 100938 280422 101494
rect 277370 78938 277606 79174
rect 277370 78618 277606 78854
rect 276146 61218 276702 61774
rect 279866 64938 280422 65494
rect 277370 42938 277606 43174
rect 277370 42618 277606 42854
rect 276146 25218 276702 25774
rect 279866 28938 280422 29494
rect 277370 6938 277606 7174
rect 277370 6618 277606 6854
rect 276146 -6662 276702 -6106
rect 279866 -7622 280422 -7066
rect 289826 704282 290382 704838
rect 289826 686898 290382 687454
rect 289826 650898 290382 651454
rect 289826 614898 290382 615454
rect 289826 578898 290382 579454
rect 289826 542898 290382 543454
rect 289826 506898 290382 507454
rect 289826 470898 290382 471454
rect 289826 434898 290382 435454
rect 289826 398898 290382 399454
rect 289826 362898 290382 363454
rect 293546 705242 294102 705798
rect 293546 690618 294102 691174
rect 293546 654618 294102 655174
rect 293546 618618 294102 619174
rect 293546 582618 294102 583174
rect 293546 546618 294102 547174
rect 293546 510618 294102 511174
rect 293546 474618 294102 475174
rect 293546 438618 294102 439174
rect 293546 402618 294102 403174
rect 293546 366618 294102 367174
rect 293546 330618 294102 331174
rect 289826 326898 290382 327454
rect 292730 327218 292966 327454
rect 292730 326898 292966 327134
rect 293546 294618 294102 295174
rect 289826 290898 290382 291454
rect 292730 291218 292966 291454
rect 292730 290898 292966 291134
rect 293546 258618 294102 259174
rect 289826 254898 290382 255454
rect 292730 255218 292966 255454
rect 292730 254898 292966 255134
rect 293546 222618 294102 223174
rect 289826 218898 290382 219454
rect 292730 219218 292966 219454
rect 292730 218898 292966 219134
rect 293546 186618 294102 187174
rect 289826 182898 290382 183454
rect 292730 183218 292966 183454
rect 292730 182898 292966 183134
rect 293546 150618 294102 151174
rect 289826 146898 290382 147454
rect 292730 147218 292966 147454
rect 292730 146898 292966 147134
rect 293546 114618 294102 115174
rect 289826 110898 290382 111454
rect 292730 111218 292966 111454
rect 292730 110898 292966 111134
rect 293546 78618 294102 79174
rect 289826 74898 290382 75454
rect 292730 75218 292966 75454
rect 292730 74898 292966 75134
rect 293546 42618 294102 43174
rect 289826 38898 290382 39454
rect 292730 39218 292966 39454
rect 292730 38898 292966 39134
rect 289826 2898 290382 3454
rect 289826 -902 290382 -346
rect 293546 6618 294102 7174
rect 293546 -1862 294102 -1306
rect 297266 706202 297822 706758
rect 297266 694338 297822 694894
rect 297266 658338 297822 658894
rect 297266 622338 297822 622894
rect 297266 586338 297822 586894
rect 297266 550338 297822 550894
rect 297266 514338 297822 514894
rect 297266 478338 297822 478894
rect 297266 442338 297822 442894
rect 297266 406338 297822 406894
rect 297266 370338 297822 370894
rect 297266 334338 297822 334894
rect 297266 298338 297822 298894
rect 297266 262338 297822 262894
rect 297266 226338 297822 226894
rect 297266 190338 297822 190894
rect 297266 154338 297822 154894
rect 297266 118338 297822 118894
rect 297266 82338 297822 82894
rect 297266 46338 297822 46894
rect 297266 10338 297822 10894
rect 297266 -2822 297822 -2266
rect 300986 707162 301542 707718
rect 300986 698058 301542 698614
rect 300986 662058 301542 662614
rect 300986 626058 301542 626614
rect 300986 590058 301542 590614
rect 300986 554058 301542 554614
rect 300986 518058 301542 518614
rect 300986 482058 301542 482614
rect 300986 446058 301542 446614
rect 300986 410058 301542 410614
rect 300986 374058 301542 374614
rect 300986 338058 301542 338614
rect 300986 302058 301542 302614
rect 300986 266058 301542 266614
rect 300986 230058 301542 230614
rect 300986 194058 301542 194614
rect 300986 158058 301542 158614
rect 300986 122058 301542 122614
rect 300986 86058 301542 86614
rect 300986 50058 301542 50614
rect 300986 14058 301542 14614
rect 300986 -3782 301542 -3226
rect 304706 708122 305262 708678
rect 304706 665778 305262 666334
rect 304706 629778 305262 630334
rect 304706 593778 305262 594334
rect 304706 557778 305262 558334
rect 304706 521778 305262 522334
rect 304706 485778 305262 486334
rect 304706 449778 305262 450334
rect 304706 413778 305262 414334
rect 304706 377778 305262 378334
rect 308426 709082 308982 709638
rect 308426 669498 308982 670054
rect 308426 633498 308982 634054
rect 308426 597498 308982 598054
rect 308426 561498 308982 562054
rect 308426 525498 308982 526054
rect 308426 489498 308982 490054
rect 308426 453498 308982 454054
rect 308426 417498 308982 418054
rect 308426 381498 308982 382054
rect 312146 710042 312702 710598
rect 312146 673218 312702 673774
rect 312146 637218 312702 637774
rect 312146 601218 312702 601774
rect 312146 565218 312702 565774
rect 312146 529218 312702 529774
rect 312146 493218 312702 493774
rect 312146 457218 312702 457774
rect 312146 421218 312702 421774
rect 312146 385218 312702 385774
rect 304706 341778 305262 342334
rect 312146 349218 312702 349774
rect 308090 330938 308326 331174
rect 308090 330618 308326 330854
rect 304706 305778 305262 306334
rect 312146 313218 312702 313774
rect 308090 294938 308326 295174
rect 308090 294618 308326 294854
rect 304706 269778 305262 270334
rect 312146 277218 312702 277774
rect 308090 258938 308326 259174
rect 308090 258618 308326 258854
rect 304706 233778 305262 234334
rect 312146 241218 312702 241774
rect 308090 222938 308326 223174
rect 308090 222618 308326 222854
rect 304706 197778 305262 198334
rect 312146 205218 312702 205774
rect 308090 186938 308326 187174
rect 308090 186618 308326 186854
rect 304706 161778 305262 162334
rect 312146 169218 312702 169774
rect 308090 150938 308326 151174
rect 308090 150618 308326 150854
rect 304706 125778 305262 126334
rect 312146 133218 312702 133774
rect 308090 114938 308326 115174
rect 308090 114618 308326 114854
rect 304706 89778 305262 90334
rect 312146 97218 312702 97774
rect 308090 78938 308326 79174
rect 308090 78618 308326 78854
rect 304706 53778 305262 54334
rect 312146 61218 312702 61774
rect 308090 42938 308326 43174
rect 308090 42618 308326 42854
rect 304706 17778 305262 18334
rect 312146 25218 312702 25774
rect 308090 6938 308326 7174
rect 308090 6618 308326 6854
rect 304706 -4742 305262 -4186
rect 312146 -6662 312702 -6106
rect 315866 711002 316422 711558
rect 315866 676938 316422 677494
rect 315866 640938 316422 641494
rect 315866 604938 316422 605494
rect 315866 568938 316422 569494
rect 315866 532938 316422 533494
rect 315866 496938 316422 497494
rect 315866 460938 316422 461494
rect 315866 424938 316422 425494
rect 315866 388938 316422 389494
rect 315866 352938 316422 353494
rect 325826 704282 326382 704838
rect 325826 686898 326382 687454
rect 325826 650898 326382 651454
rect 325826 614898 326382 615454
rect 325826 578898 326382 579454
rect 325826 542898 326382 543454
rect 325826 506898 326382 507454
rect 325826 470898 326382 471454
rect 325826 434898 326382 435454
rect 325826 398898 326382 399454
rect 325826 362898 326382 363454
rect 323450 327218 323686 327454
rect 323450 326898 323686 327134
rect 325826 326898 326382 327454
rect 315866 316938 316422 317494
rect 323450 291218 323686 291454
rect 323450 290898 323686 291134
rect 325826 290898 326382 291454
rect 315866 280938 316422 281494
rect 323450 255218 323686 255454
rect 323450 254898 323686 255134
rect 325826 254898 326382 255454
rect 315866 244938 316422 245494
rect 323450 219218 323686 219454
rect 323450 218898 323686 219134
rect 325826 218898 326382 219454
rect 315866 208938 316422 209494
rect 323450 183218 323686 183454
rect 323450 182898 323686 183134
rect 325826 182898 326382 183454
rect 315866 172938 316422 173494
rect 323450 147218 323686 147454
rect 323450 146898 323686 147134
rect 325826 146898 326382 147454
rect 315866 136938 316422 137494
rect 323450 111218 323686 111454
rect 323450 110898 323686 111134
rect 325826 110898 326382 111454
rect 315866 100938 316422 101494
rect 323450 75218 323686 75454
rect 323450 74898 323686 75134
rect 325826 74898 326382 75454
rect 315866 64938 316422 65494
rect 323450 39218 323686 39454
rect 323450 38898 323686 39134
rect 325826 38898 326382 39454
rect 315866 28938 316422 29494
rect 315866 -7622 316422 -7066
rect 325826 2898 326382 3454
rect 325826 -902 326382 -346
rect 329546 705242 330102 705798
rect 329546 690618 330102 691174
rect 329546 654618 330102 655174
rect 329546 618618 330102 619174
rect 329546 582618 330102 583174
rect 329546 546618 330102 547174
rect 329546 510618 330102 511174
rect 329546 474618 330102 475174
rect 329546 438618 330102 439174
rect 329546 402618 330102 403174
rect 329546 366618 330102 367174
rect 329546 330618 330102 331174
rect 329546 294618 330102 295174
rect 329546 258618 330102 259174
rect 329546 222618 330102 223174
rect 329546 186618 330102 187174
rect 329546 150618 330102 151174
rect 329546 114618 330102 115174
rect 329546 78618 330102 79174
rect 329546 42618 330102 43174
rect 329546 6618 330102 7174
rect 329546 -1862 330102 -1306
rect 333266 706202 333822 706758
rect 333266 694338 333822 694894
rect 333266 658338 333822 658894
rect 333266 622338 333822 622894
rect 333266 586338 333822 586894
rect 333266 550338 333822 550894
rect 333266 514338 333822 514894
rect 333266 478338 333822 478894
rect 333266 442338 333822 442894
rect 333266 406338 333822 406894
rect 333266 370338 333822 370894
rect 333266 334338 333822 334894
rect 333266 298338 333822 298894
rect 333266 262338 333822 262894
rect 333266 226338 333822 226894
rect 333266 190338 333822 190894
rect 333266 154338 333822 154894
rect 333266 118338 333822 118894
rect 333266 82338 333822 82894
rect 333266 46338 333822 46894
rect 333266 10338 333822 10894
rect 333266 -2822 333822 -2266
rect 336986 707162 337542 707718
rect 336986 698058 337542 698614
rect 336986 662058 337542 662614
rect 336986 626058 337542 626614
rect 336986 590058 337542 590614
rect 336986 554058 337542 554614
rect 336986 518058 337542 518614
rect 336986 482058 337542 482614
rect 336986 446058 337542 446614
rect 336986 410058 337542 410614
rect 336986 374058 337542 374614
rect 336986 338058 337542 338614
rect 340706 708122 341262 708678
rect 340706 665778 341262 666334
rect 340706 629778 341262 630334
rect 340706 593778 341262 594334
rect 340706 557778 341262 558334
rect 340706 521778 341262 522334
rect 340706 485778 341262 486334
rect 340706 449778 341262 450334
rect 340706 413778 341262 414334
rect 340706 377778 341262 378334
rect 340706 341778 341262 342334
rect 338810 330938 339046 331174
rect 338810 330618 339046 330854
rect 336986 302058 337542 302614
rect 340706 305778 341262 306334
rect 338810 294938 339046 295174
rect 338810 294618 339046 294854
rect 336986 266058 337542 266614
rect 340706 269778 341262 270334
rect 338810 258938 339046 259174
rect 338810 258618 339046 258854
rect 336986 230058 337542 230614
rect 340706 233778 341262 234334
rect 338810 222938 339046 223174
rect 338810 222618 339046 222854
rect 336986 194058 337542 194614
rect 340706 197778 341262 198334
rect 338810 186938 339046 187174
rect 338810 186618 339046 186854
rect 336986 158058 337542 158614
rect 340706 161778 341262 162334
rect 338810 150938 339046 151174
rect 338810 150618 339046 150854
rect 336986 122058 337542 122614
rect 340706 125778 341262 126334
rect 338810 114938 339046 115174
rect 338810 114618 339046 114854
rect 336986 86058 337542 86614
rect 340706 89778 341262 90334
rect 338810 78938 339046 79174
rect 338810 78618 339046 78854
rect 336986 50058 337542 50614
rect 340706 53778 341262 54334
rect 338810 42938 339046 43174
rect 338810 42618 339046 42854
rect 336986 14058 337542 14614
rect 340706 17778 341262 18334
rect 338810 6938 339046 7174
rect 338810 6618 339046 6854
rect 336986 -3782 337542 -3226
rect 340706 -4742 341262 -4186
rect 344426 709082 344982 709638
rect 344426 669498 344982 670054
rect 344426 633498 344982 634054
rect 344426 597498 344982 598054
rect 344426 561498 344982 562054
rect 344426 525498 344982 526054
rect 344426 489498 344982 490054
rect 344426 453498 344982 454054
rect 344426 417498 344982 418054
rect 344426 381498 344982 382054
rect 344426 345498 344982 346054
rect 344426 309498 344982 310054
rect 344426 273498 344982 274054
rect 344426 237498 344982 238054
rect 344426 201498 344982 202054
rect 344426 165498 344982 166054
rect 344426 129498 344982 130054
rect 344426 93498 344982 94054
rect 344426 57498 344982 58054
rect 344426 21498 344982 22054
rect 344426 -5702 344982 -5146
rect 348146 710042 348702 710598
rect 348146 673218 348702 673774
rect 348146 637218 348702 637774
rect 348146 601218 348702 601774
rect 348146 565218 348702 565774
rect 348146 529218 348702 529774
rect 348146 493218 348702 493774
rect 348146 457218 348702 457774
rect 348146 421218 348702 421774
rect 348146 385218 348702 385774
rect 348146 349218 348702 349774
rect 348146 313218 348702 313774
rect 348146 277218 348702 277774
rect 348146 241218 348702 241774
rect 348146 205218 348702 205774
rect 348146 169218 348702 169774
rect 348146 133218 348702 133774
rect 348146 97218 348702 97774
rect 348146 61218 348702 61774
rect 348146 25218 348702 25774
rect 348146 -6662 348702 -6106
rect 351866 711002 352422 711558
rect 351866 676938 352422 677494
rect 351866 640938 352422 641494
rect 351866 604938 352422 605494
rect 351866 568938 352422 569494
rect 351866 532938 352422 533494
rect 351866 496938 352422 497494
rect 351866 460938 352422 461494
rect 351866 424938 352422 425494
rect 351866 388938 352422 389494
rect 351866 352938 352422 353494
rect 361826 704282 362382 704838
rect 361826 686898 362382 687454
rect 361826 650898 362382 651454
rect 361826 614898 362382 615454
rect 361826 578898 362382 579454
rect 361826 542898 362382 543454
rect 361826 506898 362382 507454
rect 361826 470898 362382 471454
rect 361826 434898 362382 435454
rect 361826 398898 362382 399454
rect 361826 362898 362382 363454
rect 354170 327218 354406 327454
rect 354170 326898 354406 327134
rect 361826 326898 362382 327454
rect 351866 316938 352422 317494
rect 354170 291218 354406 291454
rect 354170 290898 354406 291134
rect 361826 290898 362382 291454
rect 351866 280938 352422 281494
rect 354170 255218 354406 255454
rect 354170 254898 354406 255134
rect 361826 254898 362382 255454
rect 351866 244938 352422 245494
rect 354170 219218 354406 219454
rect 354170 218898 354406 219134
rect 361826 218898 362382 219454
rect 351866 208938 352422 209494
rect 354170 183218 354406 183454
rect 354170 182898 354406 183134
rect 361826 182898 362382 183454
rect 351866 172938 352422 173494
rect 354170 147218 354406 147454
rect 354170 146898 354406 147134
rect 361826 146898 362382 147454
rect 351866 136938 352422 137494
rect 354170 111218 354406 111454
rect 354170 110898 354406 111134
rect 361826 110898 362382 111454
rect 351866 100938 352422 101494
rect 354170 75218 354406 75454
rect 354170 74898 354406 75134
rect 361826 74898 362382 75454
rect 351866 64938 352422 65494
rect 354170 39218 354406 39454
rect 354170 38898 354406 39134
rect 361826 38898 362382 39454
rect 351866 28938 352422 29494
rect 351866 -7622 352422 -7066
rect 361826 2898 362382 3454
rect 361826 -902 362382 -346
rect 365546 705242 366102 705798
rect 365546 690618 366102 691174
rect 365546 654618 366102 655174
rect 365546 618618 366102 619174
rect 365546 582618 366102 583174
rect 365546 546618 366102 547174
rect 365546 510618 366102 511174
rect 365546 474618 366102 475174
rect 365546 438618 366102 439174
rect 365546 402618 366102 403174
rect 365546 366618 366102 367174
rect 369266 706202 369822 706758
rect 369266 694338 369822 694894
rect 369266 658338 369822 658894
rect 369266 622338 369822 622894
rect 369266 586338 369822 586894
rect 369266 550338 369822 550894
rect 369266 514338 369822 514894
rect 369266 478338 369822 478894
rect 369266 442338 369822 442894
rect 369266 406338 369822 406894
rect 369266 370338 369822 370894
rect 372986 707162 373542 707718
rect 372986 698058 373542 698614
rect 372986 662058 373542 662614
rect 372986 626058 373542 626614
rect 372986 590058 373542 590614
rect 372986 554058 373542 554614
rect 372986 518058 373542 518614
rect 372986 482058 373542 482614
rect 372986 446058 373542 446614
rect 372986 410058 373542 410614
rect 372986 374058 373542 374614
rect 372986 338058 373542 338614
rect 365546 330618 366102 331174
rect 369530 330938 369766 331174
rect 369530 330618 369766 330854
rect 372986 302058 373542 302614
rect 365546 294618 366102 295174
rect 369530 294938 369766 295174
rect 369530 294618 369766 294854
rect 372986 266058 373542 266614
rect 365546 258618 366102 259174
rect 369530 258938 369766 259174
rect 369530 258618 369766 258854
rect 372986 230058 373542 230614
rect 365546 222618 366102 223174
rect 369530 222938 369766 223174
rect 369530 222618 369766 222854
rect 372986 194058 373542 194614
rect 365546 186618 366102 187174
rect 369530 186938 369766 187174
rect 369530 186618 369766 186854
rect 372986 158058 373542 158614
rect 365546 150618 366102 151174
rect 369530 150938 369766 151174
rect 369530 150618 369766 150854
rect 372986 122058 373542 122614
rect 365546 114618 366102 115174
rect 369530 114938 369766 115174
rect 369530 114618 369766 114854
rect 372986 86058 373542 86614
rect 365546 78618 366102 79174
rect 369530 78938 369766 79174
rect 369530 78618 369766 78854
rect 372986 50058 373542 50614
rect 365546 42618 366102 43174
rect 369530 42938 369766 43174
rect 369530 42618 369766 42854
rect 372986 14058 373542 14614
rect 365546 6618 366102 7174
rect 369530 6938 369766 7174
rect 369530 6618 369766 6854
rect 365546 -1862 366102 -1306
rect 372986 -3782 373542 -3226
rect 376706 708122 377262 708678
rect 376706 665778 377262 666334
rect 376706 629778 377262 630334
rect 376706 593778 377262 594334
rect 376706 557778 377262 558334
rect 376706 521778 377262 522334
rect 376706 485778 377262 486334
rect 376706 449778 377262 450334
rect 376706 413778 377262 414334
rect 376706 377778 377262 378334
rect 376706 341778 377262 342334
rect 376706 305778 377262 306334
rect 376706 269778 377262 270334
rect 376706 233778 377262 234334
rect 376706 197778 377262 198334
rect 376706 161778 377262 162334
rect 376706 125778 377262 126334
rect 376706 89778 377262 90334
rect 376706 53778 377262 54334
rect 376706 17778 377262 18334
rect 376706 -4742 377262 -4186
rect 380426 709082 380982 709638
rect 380426 669498 380982 670054
rect 380426 633498 380982 634054
rect 380426 597498 380982 598054
rect 380426 561498 380982 562054
rect 380426 525498 380982 526054
rect 380426 489498 380982 490054
rect 380426 453498 380982 454054
rect 380426 417498 380982 418054
rect 380426 381498 380982 382054
rect 380426 345498 380982 346054
rect 380426 309498 380982 310054
rect 380426 273498 380982 274054
rect 380426 237498 380982 238054
rect 380426 201498 380982 202054
rect 380426 165498 380982 166054
rect 380426 129498 380982 130054
rect 380426 93498 380982 94054
rect 380426 57498 380982 58054
rect 380426 21498 380982 22054
rect 380426 -5702 380982 -5146
rect 384146 710042 384702 710598
rect 384146 673218 384702 673774
rect 384146 637218 384702 637774
rect 384146 601218 384702 601774
rect 384146 565218 384702 565774
rect 384146 529218 384702 529774
rect 384146 493218 384702 493774
rect 384146 457218 384702 457774
rect 384146 421218 384702 421774
rect 384146 385218 384702 385774
rect 384146 349218 384702 349774
rect 387866 711002 388422 711558
rect 387866 676938 388422 677494
rect 387866 640938 388422 641494
rect 387866 604938 388422 605494
rect 387866 568938 388422 569494
rect 387866 532938 388422 533494
rect 387866 496938 388422 497494
rect 387866 460938 388422 461494
rect 387866 424938 388422 425494
rect 387866 388938 388422 389494
rect 387866 352938 388422 353494
rect 384890 327218 385126 327454
rect 384890 326898 385126 327134
rect 384146 313218 384702 313774
rect 387866 316938 388422 317494
rect 384890 291218 385126 291454
rect 384890 290898 385126 291134
rect 384146 277218 384702 277774
rect 387866 280938 388422 281494
rect 384890 255218 385126 255454
rect 384890 254898 385126 255134
rect 384146 241218 384702 241774
rect 387866 244938 388422 245494
rect 384890 219218 385126 219454
rect 384890 218898 385126 219134
rect 384146 205218 384702 205774
rect 387866 208938 388422 209494
rect 384890 183218 385126 183454
rect 384890 182898 385126 183134
rect 384146 169218 384702 169774
rect 387866 172938 388422 173494
rect 384890 147218 385126 147454
rect 384890 146898 385126 147134
rect 384146 133218 384702 133774
rect 387866 136938 388422 137494
rect 384890 111218 385126 111454
rect 384890 110898 385126 111134
rect 384146 97218 384702 97774
rect 387866 100938 388422 101494
rect 384890 75218 385126 75454
rect 384890 74898 385126 75134
rect 384146 61218 384702 61774
rect 387866 64938 388422 65494
rect 384890 39218 385126 39454
rect 384890 38898 385126 39134
rect 384146 25218 384702 25774
rect 384146 -6662 384702 -6106
rect 387866 28938 388422 29494
rect 387866 -7622 388422 -7066
rect 397826 704282 398382 704838
rect 397826 686898 398382 687454
rect 397826 650898 398382 651454
rect 397826 614898 398382 615454
rect 397826 578898 398382 579454
rect 397826 542898 398382 543454
rect 397826 506898 398382 507454
rect 397826 470898 398382 471454
rect 397826 434898 398382 435454
rect 397826 398898 398382 399454
rect 397826 362898 398382 363454
rect 401546 705242 402102 705798
rect 401546 690618 402102 691174
rect 401546 654618 402102 655174
rect 401546 618618 402102 619174
rect 401546 582618 402102 583174
rect 401546 546618 402102 547174
rect 401546 510618 402102 511174
rect 401546 474618 402102 475174
rect 401546 438618 402102 439174
rect 401546 402618 402102 403174
rect 401546 366618 402102 367174
rect 400250 330938 400486 331174
rect 400250 330618 400486 330854
rect 401546 330618 402102 331174
rect 397826 326898 398382 327454
rect 400250 294938 400486 295174
rect 400250 294618 400486 294854
rect 401546 294618 402102 295174
rect 397826 290898 398382 291454
rect 400250 258938 400486 259174
rect 400250 258618 400486 258854
rect 401546 258618 402102 259174
rect 397826 254898 398382 255454
rect 400250 222938 400486 223174
rect 400250 222618 400486 222854
rect 401546 222618 402102 223174
rect 397826 218898 398382 219454
rect 400250 186938 400486 187174
rect 400250 186618 400486 186854
rect 401546 186618 402102 187174
rect 397826 182898 398382 183454
rect 400250 150938 400486 151174
rect 400250 150618 400486 150854
rect 401546 150618 402102 151174
rect 397826 146898 398382 147454
rect 400250 114938 400486 115174
rect 400250 114618 400486 114854
rect 401546 114618 402102 115174
rect 397826 110898 398382 111454
rect 400250 78938 400486 79174
rect 400250 78618 400486 78854
rect 401546 78618 402102 79174
rect 397826 74898 398382 75454
rect 400250 42938 400486 43174
rect 400250 42618 400486 42854
rect 401546 42618 402102 43174
rect 397826 38898 398382 39454
rect 400250 6938 400486 7174
rect 400250 6618 400486 6854
rect 401546 6618 402102 7174
rect 397826 2898 398382 3454
rect 397826 -902 398382 -346
rect 401546 -1862 402102 -1306
rect 405266 706202 405822 706758
rect 405266 694338 405822 694894
rect 405266 658338 405822 658894
rect 405266 622338 405822 622894
rect 405266 586338 405822 586894
rect 405266 550338 405822 550894
rect 405266 514338 405822 514894
rect 405266 478338 405822 478894
rect 405266 442338 405822 442894
rect 405266 406338 405822 406894
rect 405266 370338 405822 370894
rect 405266 334338 405822 334894
rect 405266 298338 405822 298894
rect 405266 262338 405822 262894
rect 405266 226338 405822 226894
rect 405266 190338 405822 190894
rect 405266 154338 405822 154894
rect 405266 118338 405822 118894
rect 405266 82338 405822 82894
rect 405266 46338 405822 46894
rect 405266 10338 405822 10894
rect 405266 -2822 405822 -2266
rect 408986 707162 409542 707718
rect 408986 698058 409542 698614
rect 408986 662058 409542 662614
rect 408986 626058 409542 626614
rect 408986 590058 409542 590614
rect 408986 554058 409542 554614
rect 408986 518058 409542 518614
rect 408986 482058 409542 482614
rect 408986 446058 409542 446614
rect 408986 410058 409542 410614
rect 408986 374058 409542 374614
rect 408986 338058 409542 338614
rect 408986 302058 409542 302614
rect 408986 266058 409542 266614
rect 408986 230058 409542 230614
rect 408986 194058 409542 194614
rect 408986 158058 409542 158614
rect 408986 122058 409542 122614
rect 408986 86058 409542 86614
rect 408986 50058 409542 50614
rect 408986 14058 409542 14614
rect 408986 -3782 409542 -3226
rect 412706 708122 413262 708678
rect 412706 665778 413262 666334
rect 412706 629778 413262 630334
rect 412706 593778 413262 594334
rect 412706 557778 413262 558334
rect 412706 521778 413262 522334
rect 412706 485778 413262 486334
rect 412706 449778 413262 450334
rect 412706 413778 413262 414334
rect 412706 377778 413262 378334
rect 412706 341778 413262 342334
rect 416426 709082 416982 709638
rect 416426 669498 416982 670054
rect 416426 633498 416982 634054
rect 416426 597498 416982 598054
rect 416426 561498 416982 562054
rect 416426 525498 416982 526054
rect 416426 489498 416982 490054
rect 416426 453498 416982 454054
rect 416426 417498 416982 418054
rect 416426 381498 416982 382054
rect 416426 345498 416982 346054
rect 415610 327218 415846 327454
rect 415610 326898 415846 327134
rect 412706 305778 413262 306334
rect 416426 309498 416982 310054
rect 415610 291218 415846 291454
rect 415610 290898 415846 291134
rect 412706 269778 413262 270334
rect 416426 273498 416982 274054
rect 415610 255218 415846 255454
rect 415610 254898 415846 255134
rect 412706 233778 413262 234334
rect 416426 237498 416982 238054
rect 415610 219218 415846 219454
rect 415610 218898 415846 219134
rect 412706 197778 413262 198334
rect 416426 201498 416982 202054
rect 415610 183218 415846 183454
rect 415610 182898 415846 183134
rect 412706 161778 413262 162334
rect 416426 165498 416982 166054
rect 415610 147218 415846 147454
rect 415610 146898 415846 147134
rect 412706 125778 413262 126334
rect 416426 129498 416982 130054
rect 415610 111218 415846 111454
rect 415610 110898 415846 111134
rect 412706 89778 413262 90334
rect 416426 93498 416982 94054
rect 415610 75218 415846 75454
rect 415610 74898 415846 75134
rect 412706 53778 413262 54334
rect 416426 57498 416982 58054
rect 415610 39218 415846 39454
rect 415610 38898 415846 39134
rect 412706 17778 413262 18334
rect 412706 -4742 413262 -4186
rect 416426 21498 416982 22054
rect 416426 -5702 416982 -5146
rect 420146 710042 420702 710598
rect 420146 673218 420702 673774
rect 420146 637218 420702 637774
rect 420146 601218 420702 601774
rect 420146 565218 420702 565774
rect 420146 529218 420702 529774
rect 420146 493218 420702 493774
rect 420146 457218 420702 457774
rect 420146 421218 420702 421774
rect 420146 385218 420702 385774
rect 420146 349218 420702 349774
rect 420146 313218 420702 313774
rect 420146 277218 420702 277774
rect 420146 241218 420702 241774
rect 420146 205218 420702 205774
rect 420146 169218 420702 169774
rect 420146 133218 420702 133774
rect 420146 97218 420702 97774
rect 420146 61218 420702 61774
rect 420146 25218 420702 25774
rect 420146 -6662 420702 -6106
rect 423866 711002 424422 711558
rect 423866 676938 424422 677494
rect 423866 640938 424422 641494
rect 423866 604938 424422 605494
rect 423866 568938 424422 569494
rect 423866 532938 424422 533494
rect 423866 496938 424422 497494
rect 423866 460938 424422 461494
rect 423866 424938 424422 425494
rect 423866 388938 424422 389494
rect 423866 352938 424422 353494
rect 433826 704282 434382 704838
rect 433826 686898 434382 687454
rect 433826 650898 434382 651454
rect 433826 614898 434382 615454
rect 433826 578898 434382 579454
rect 433826 542898 434382 543454
rect 433826 506898 434382 507454
rect 433826 470898 434382 471454
rect 433826 434898 434382 435454
rect 433826 398898 434382 399454
rect 433826 362898 434382 363454
rect 430970 330938 431206 331174
rect 430970 330618 431206 330854
rect 423866 316938 424422 317494
rect 433826 326898 434382 327454
rect 430970 294938 431206 295174
rect 430970 294618 431206 294854
rect 423866 280938 424422 281494
rect 433826 290898 434382 291454
rect 430970 258938 431206 259174
rect 430970 258618 431206 258854
rect 423866 244938 424422 245494
rect 433826 254898 434382 255454
rect 430970 222938 431206 223174
rect 430970 222618 431206 222854
rect 423866 208938 424422 209494
rect 433826 218898 434382 219454
rect 430970 186938 431206 187174
rect 430970 186618 431206 186854
rect 423866 172938 424422 173494
rect 433826 182898 434382 183454
rect 430970 150938 431206 151174
rect 430970 150618 431206 150854
rect 423866 136938 424422 137494
rect 433826 146898 434382 147454
rect 430970 114938 431206 115174
rect 430970 114618 431206 114854
rect 423866 100938 424422 101494
rect 433826 110898 434382 111454
rect 430970 78938 431206 79174
rect 430970 78618 431206 78854
rect 423866 64938 424422 65494
rect 433826 74898 434382 75454
rect 430970 42938 431206 43174
rect 430970 42618 431206 42854
rect 423866 28938 424422 29494
rect 433826 38898 434382 39454
rect 430970 6938 431206 7174
rect 430970 6618 431206 6854
rect 423866 -7622 424422 -7066
rect 433826 2898 434382 3454
rect 433826 -902 434382 -346
rect 437546 705242 438102 705798
rect 437546 690618 438102 691174
rect 437546 654618 438102 655174
rect 437546 618618 438102 619174
rect 437546 582618 438102 583174
rect 437546 546618 438102 547174
rect 437546 510618 438102 511174
rect 437546 474618 438102 475174
rect 437546 438618 438102 439174
rect 437546 402618 438102 403174
rect 437546 366618 438102 367174
rect 437546 330618 438102 331174
rect 437546 294618 438102 295174
rect 437546 258618 438102 259174
rect 437546 222618 438102 223174
rect 437546 186618 438102 187174
rect 437546 150618 438102 151174
rect 437546 114618 438102 115174
rect 437546 78618 438102 79174
rect 437546 42618 438102 43174
rect 437546 6618 438102 7174
rect 437546 -1862 438102 -1306
rect 441266 706202 441822 706758
rect 441266 694338 441822 694894
rect 441266 658338 441822 658894
rect 441266 622338 441822 622894
rect 441266 586338 441822 586894
rect 441266 550338 441822 550894
rect 441266 514338 441822 514894
rect 441266 478338 441822 478894
rect 441266 442338 441822 442894
rect 441266 406338 441822 406894
rect 441266 370338 441822 370894
rect 441266 334338 441822 334894
rect 441266 298338 441822 298894
rect 441266 262338 441822 262894
rect 441266 226338 441822 226894
rect 441266 190338 441822 190894
rect 441266 154338 441822 154894
rect 441266 118338 441822 118894
rect 441266 82338 441822 82894
rect 441266 46338 441822 46894
rect 441266 10338 441822 10894
rect 441266 -2822 441822 -2266
rect 444986 707162 445542 707718
rect 444986 698058 445542 698614
rect 444986 662058 445542 662614
rect 444986 626058 445542 626614
rect 444986 590058 445542 590614
rect 444986 554058 445542 554614
rect 444986 518058 445542 518614
rect 444986 482058 445542 482614
rect 444986 446058 445542 446614
rect 444986 410058 445542 410614
rect 444986 374058 445542 374614
rect 444986 338058 445542 338614
rect 448706 708122 449262 708678
rect 448706 665778 449262 666334
rect 448706 629778 449262 630334
rect 448706 593778 449262 594334
rect 448706 557778 449262 558334
rect 448706 521778 449262 522334
rect 448706 485778 449262 486334
rect 448706 449778 449262 450334
rect 448706 413778 449262 414334
rect 448706 377778 449262 378334
rect 448706 341778 449262 342334
rect 446330 327218 446566 327454
rect 446330 326898 446566 327134
rect 444986 302058 445542 302614
rect 448706 305778 449262 306334
rect 446330 291218 446566 291454
rect 446330 290898 446566 291134
rect 444986 266058 445542 266614
rect 448706 269778 449262 270334
rect 446330 255218 446566 255454
rect 446330 254898 446566 255134
rect 444986 230058 445542 230614
rect 448706 233778 449262 234334
rect 446330 219218 446566 219454
rect 446330 218898 446566 219134
rect 444986 194058 445542 194614
rect 448706 197778 449262 198334
rect 446330 183218 446566 183454
rect 446330 182898 446566 183134
rect 444986 158058 445542 158614
rect 448706 161778 449262 162334
rect 446330 147218 446566 147454
rect 446330 146898 446566 147134
rect 444986 122058 445542 122614
rect 448706 125778 449262 126334
rect 446330 111218 446566 111454
rect 446330 110898 446566 111134
rect 444986 86058 445542 86614
rect 448706 89778 449262 90334
rect 446330 75218 446566 75454
rect 446330 74898 446566 75134
rect 444986 50058 445542 50614
rect 448706 53778 449262 54334
rect 446330 39218 446566 39454
rect 446330 38898 446566 39134
rect 444986 14058 445542 14614
rect 444986 -3782 445542 -3226
rect 448706 17778 449262 18334
rect 448706 -4742 449262 -4186
rect 452426 709082 452982 709638
rect 452426 669498 452982 670054
rect 452426 633498 452982 634054
rect 452426 597498 452982 598054
rect 452426 561498 452982 562054
rect 452426 525498 452982 526054
rect 452426 489498 452982 490054
rect 452426 453498 452982 454054
rect 452426 417498 452982 418054
rect 452426 381498 452982 382054
rect 452426 345498 452982 346054
rect 452426 309498 452982 310054
rect 452426 273498 452982 274054
rect 452426 237498 452982 238054
rect 452426 201498 452982 202054
rect 452426 165498 452982 166054
rect 452426 129498 452982 130054
rect 452426 93498 452982 94054
rect 452426 57498 452982 58054
rect 452426 21498 452982 22054
rect 452426 -5702 452982 -5146
rect 456146 710042 456702 710598
rect 456146 673218 456702 673774
rect 456146 637218 456702 637774
rect 456146 601218 456702 601774
rect 456146 565218 456702 565774
rect 456146 529218 456702 529774
rect 456146 493218 456702 493774
rect 456146 457218 456702 457774
rect 456146 421218 456702 421774
rect 456146 385218 456702 385774
rect 456146 349218 456702 349774
rect 456146 313218 456702 313774
rect 456146 277218 456702 277774
rect 456146 241218 456702 241774
rect 456146 205218 456702 205774
rect 456146 169218 456702 169774
rect 456146 133218 456702 133774
rect 456146 97218 456702 97774
rect 456146 61218 456702 61774
rect 456146 25218 456702 25774
rect 456146 -6662 456702 -6106
rect 459866 711002 460422 711558
rect 459866 676938 460422 677494
rect 459866 640938 460422 641494
rect 459866 604938 460422 605494
rect 459866 568938 460422 569494
rect 459866 532938 460422 533494
rect 459866 496938 460422 497494
rect 459866 460938 460422 461494
rect 459866 424938 460422 425494
rect 459866 388938 460422 389494
rect 459866 352938 460422 353494
rect 469826 704282 470382 704838
rect 469826 686898 470382 687454
rect 469826 650898 470382 651454
rect 469826 614898 470382 615454
rect 469826 578898 470382 579454
rect 469826 542898 470382 543454
rect 469826 506898 470382 507454
rect 469826 470898 470382 471454
rect 469826 434898 470382 435454
rect 469826 398898 470382 399454
rect 469826 362898 470382 363454
rect 461690 330938 461926 331174
rect 461690 330618 461926 330854
rect 459866 316938 460422 317494
rect 469826 326898 470382 327454
rect 461690 294938 461926 295174
rect 461690 294618 461926 294854
rect 459866 280938 460422 281494
rect 469826 290898 470382 291454
rect 461690 258938 461926 259174
rect 461690 258618 461926 258854
rect 459866 244938 460422 245494
rect 469826 254898 470382 255454
rect 461690 222938 461926 223174
rect 461690 222618 461926 222854
rect 459866 208938 460422 209494
rect 469826 218898 470382 219454
rect 461690 186938 461926 187174
rect 461690 186618 461926 186854
rect 459866 172938 460422 173494
rect 469826 182898 470382 183454
rect 461690 150938 461926 151174
rect 461690 150618 461926 150854
rect 459866 136938 460422 137494
rect 469826 146898 470382 147454
rect 461690 114938 461926 115174
rect 461690 114618 461926 114854
rect 459866 100938 460422 101494
rect 469826 110898 470382 111454
rect 461690 78938 461926 79174
rect 461690 78618 461926 78854
rect 459866 64938 460422 65494
rect 469826 74898 470382 75454
rect 461690 42938 461926 43174
rect 461690 42618 461926 42854
rect 459866 28938 460422 29494
rect 469826 38898 470382 39454
rect 461690 6938 461926 7174
rect 461690 6618 461926 6854
rect 459866 -7622 460422 -7066
rect 469826 2898 470382 3454
rect 469826 -902 470382 -346
rect 473546 705242 474102 705798
rect 473546 690618 474102 691174
rect 473546 654618 474102 655174
rect 473546 618618 474102 619174
rect 473546 582618 474102 583174
rect 473546 546618 474102 547174
rect 473546 510618 474102 511174
rect 473546 474618 474102 475174
rect 473546 438618 474102 439174
rect 473546 402618 474102 403174
rect 473546 366618 474102 367174
rect 477266 706202 477822 706758
rect 477266 694338 477822 694894
rect 477266 658338 477822 658894
rect 477266 622338 477822 622894
rect 477266 586338 477822 586894
rect 477266 550338 477822 550894
rect 477266 514338 477822 514894
rect 477266 478338 477822 478894
rect 477266 442338 477822 442894
rect 477266 406338 477822 406894
rect 477266 370338 477822 370894
rect 480986 707162 481542 707718
rect 480986 698058 481542 698614
rect 480986 662058 481542 662614
rect 480986 626058 481542 626614
rect 480986 590058 481542 590614
rect 480986 554058 481542 554614
rect 480986 518058 481542 518614
rect 480986 482058 481542 482614
rect 480986 446058 481542 446614
rect 480986 410058 481542 410614
rect 480986 374058 481542 374614
rect 473546 330618 474102 331174
rect 480986 338058 481542 338614
rect 477050 327218 477286 327454
rect 477050 326898 477286 327134
rect 473546 294618 474102 295174
rect 480986 302058 481542 302614
rect 477050 291218 477286 291454
rect 477050 290898 477286 291134
rect 473546 258618 474102 259174
rect 480986 266058 481542 266614
rect 477050 255218 477286 255454
rect 477050 254898 477286 255134
rect 473546 222618 474102 223174
rect 480986 230058 481542 230614
rect 477050 219218 477286 219454
rect 477050 218898 477286 219134
rect 473546 186618 474102 187174
rect 480986 194058 481542 194614
rect 477050 183218 477286 183454
rect 477050 182898 477286 183134
rect 473546 150618 474102 151174
rect 480986 158058 481542 158614
rect 477050 147218 477286 147454
rect 477050 146898 477286 147134
rect 473546 114618 474102 115174
rect 480986 122058 481542 122614
rect 477050 111218 477286 111454
rect 477050 110898 477286 111134
rect 473546 78618 474102 79174
rect 480986 86058 481542 86614
rect 477050 75218 477286 75454
rect 477050 74898 477286 75134
rect 473546 42618 474102 43174
rect 480986 50058 481542 50614
rect 477050 39218 477286 39454
rect 477050 38898 477286 39134
rect 473546 6618 474102 7174
rect 473546 -1862 474102 -1306
rect 480986 14058 481542 14614
rect 480986 -3782 481542 -3226
rect 484706 708122 485262 708678
rect 484706 665778 485262 666334
rect 484706 629778 485262 630334
rect 484706 593778 485262 594334
rect 484706 557778 485262 558334
rect 484706 521778 485262 522334
rect 484706 485778 485262 486334
rect 484706 449778 485262 450334
rect 484706 413778 485262 414334
rect 484706 377778 485262 378334
rect 484706 341778 485262 342334
rect 484706 305778 485262 306334
rect 484706 269778 485262 270334
rect 484706 233778 485262 234334
rect 484706 197778 485262 198334
rect 484706 161778 485262 162334
rect 484706 125778 485262 126334
rect 484706 89778 485262 90334
rect 484706 53778 485262 54334
rect 484706 17778 485262 18334
rect 484706 -4742 485262 -4186
rect 488426 709082 488982 709638
rect 488426 669498 488982 670054
rect 488426 633498 488982 634054
rect 488426 597498 488982 598054
rect 488426 561498 488982 562054
rect 488426 525498 488982 526054
rect 488426 489498 488982 490054
rect 488426 453498 488982 454054
rect 488426 417498 488982 418054
rect 488426 381498 488982 382054
rect 492146 710042 492702 710598
rect 492146 673218 492702 673774
rect 492146 637218 492702 637774
rect 492146 601218 492702 601774
rect 492146 565218 492702 565774
rect 492146 529218 492702 529774
rect 492146 493218 492702 493774
rect 492146 457218 492702 457774
rect 492146 421218 492702 421774
rect 492146 385218 492702 385774
rect 495866 711002 496422 711558
rect 495866 676938 496422 677494
rect 495866 640938 496422 641494
rect 495866 604938 496422 605494
rect 495866 568938 496422 569494
rect 495866 532938 496422 533494
rect 495866 496938 496422 497494
rect 495866 460938 496422 461494
rect 495866 424938 496422 425494
rect 495866 388938 496422 389494
rect 488426 345498 488982 346054
rect 495866 352938 496422 353494
rect 492410 330938 492646 331174
rect 492410 330618 492646 330854
rect 488426 309498 488982 310054
rect 495866 316938 496422 317494
rect 492410 294938 492646 295174
rect 492410 294618 492646 294854
rect 488426 273498 488982 274054
rect 495866 280938 496422 281494
rect 492410 258938 492646 259174
rect 492410 258618 492646 258854
rect 488426 237498 488982 238054
rect 495866 244938 496422 245494
rect 492410 222938 492646 223174
rect 492410 222618 492646 222854
rect 488426 201498 488982 202054
rect 495866 208938 496422 209494
rect 492410 186938 492646 187174
rect 492410 186618 492646 186854
rect 488426 165498 488982 166054
rect 495866 172938 496422 173494
rect 492410 150938 492646 151174
rect 492410 150618 492646 150854
rect 488426 129498 488982 130054
rect 495866 136938 496422 137494
rect 492410 114938 492646 115174
rect 492410 114618 492646 114854
rect 488426 93498 488982 94054
rect 495866 100938 496422 101494
rect 492410 78938 492646 79174
rect 492410 78618 492646 78854
rect 488426 57498 488982 58054
rect 495866 64938 496422 65494
rect 492410 42938 492646 43174
rect 492410 42618 492646 42854
rect 488426 21498 488982 22054
rect 495866 28938 496422 29494
rect 492410 6938 492646 7174
rect 492410 6618 492646 6854
rect 488426 -5702 488982 -5146
rect 495866 -7622 496422 -7066
rect 505826 704282 506382 704838
rect 505826 686898 506382 687454
rect 505826 650898 506382 651454
rect 505826 614898 506382 615454
rect 505826 578898 506382 579454
rect 505826 542898 506382 543454
rect 505826 506898 506382 507454
rect 505826 470898 506382 471454
rect 505826 434898 506382 435454
rect 505826 398898 506382 399454
rect 505826 362898 506382 363454
rect 509546 705242 510102 705798
rect 509546 690618 510102 691174
rect 509546 654618 510102 655174
rect 509546 618618 510102 619174
rect 509546 582618 510102 583174
rect 509546 546618 510102 547174
rect 509546 510618 510102 511174
rect 509546 474618 510102 475174
rect 509546 438618 510102 439174
rect 509546 402618 510102 403174
rect 509546 366618 510102 367174
rect 509546 330618 510102 331174
rect 505826 326898 506382 327454
rect 507770 327218 508006 327454
rect 507770 326898 508006 327134
rect 509546 294618 510102 295174
rect 505826 290898 506382 291454
rect 507770 291218 508006 291454
rect 507770 290898 508006 291134
rect 509546 258618 510102 259174
rect 505826 254898 506382 255454
rect 507770 255218 508006 255454
rect 507770 254898 508006 255134
rect 509546 222618 510102 223174
rect 505826 218898 506382 219454
rect 507770 219218 508006 219454
rect 507770 218898 508006 219134
rect 509546 186618 510102 187174
rect 505826 182898 506382 183454
rect 507770 183218 508006 183454
rect 507770 182898 508006 183134
rect 509546 150618 510102 151174
rect 505826 146898 506382 147454
rect 507770 147218 508006 147454
rect 507770 146898 508006 147134
rect 509546 114618 510102 115174
rect 505826 110898 506382 111454
rect 507770 111218 508006 111454
rect 507770 110898 508006 111134
rect 509546 78618 510102 79174
rect 505826 74898 506382 75454
rect 507770 75218 508006 75454
rect 507770 74898 508006 75134
rect 509546 42618 510102 43174
rect 505826 38898 506382 39454
rect 507770 39218 508006 39454
rect 507770 38898 508006 39134
rect 505826 2898 506382 3454
rect 505826 -902 506382 -346
rect 509546 6618 510102 7174
rect 509546 -1862 510102 -1306
rect 513266 706202 513822 706758
rect 513266 694338 513822 694894
rect 513266 658338 513822 658894
rect 513266 622338 513822 622894
rect 513266 586338 513822 586894
rect 513266 550338 513822 550894
rect 513266 514338 513822 514894
rect 513266 478338 513822 478894
rect 513266 442338 513822 442894
rect 513266 406338 513822 406894
rect 513266 370338 513822 370894
rect 513266 334338 513822 334894
rect 513266 298338 513822 298894
rect 513266 262338 513822 262894
rect 513266 226338 513822 226894
rect 513266 190338 513822 190894
rect 513266 154338 513822 154894
rect 513266 118338 513822 118894
rect 513266 82338 513822 82894
rect 513266 46338 513822 46894
rect 513266 10338 513822 10894
rect 513266 -2822 513822 -2266
rect 516986 707162 517542 707718
rect 516986 698058 517542 698614
rect 516986 662058 517542 662614
rect 516986 626058 517542 626614
rect 516986 590058 517542 590614
rect 516986 554058 517542 554614
rect 516986 518058 517542 518614
rect 516986 482058 517542 482614
rect 516986 446058 517542 446614
rect 516986 410058 517542 410614
rect 516986 374058 517542 374614
rect 516986 338058 517542 338614
rect 516986 302058 517542 302614
rect 516986 266058 517542 266614
rect 516986 230058 517542 230614
rect 516986 194058 517542 194614
rect 516986 158058 517542 158614
rect 516986 122058 517542 122614
rect 516986 86058 517542 86614
rect 516986 50058 517542 50614
rect 516986 14058 517542 14614
rect 516986 -3782 517542 -3226
rect 520706 708122 521262 708678
rect 520706 665778 521262 666334
rect 520706 629778 521262 630334
rect 520706 593778 521262 594334
rect 520706 557778 521262 558334
rect 520706 521778 521262 522334
rect 520706 485778 521262 486334
rect 520706 449778 521262 450334
rect 520706 413778 521262 414334
rect 520706 377778 521262 378334
rect 520706 341778 521262 342334
rect 524426 709082 524982 709638
rect 524426 669498 524982 670054
rect 524426 633498 524982 634054
rect 524426 597498 524982 598054
rect 524426 561498 524982 562054
rect 524426 525498 524982 526054
rect 524426 489498 524982 490054
rect 524426 453498 524982 454054
rect 524426 417498 524982 418054
rect 524426 381498 524982 382054
rect 524426 345498 524982 346054
rect 523130 330938 523366 331174
rect 523130 330618 523366 330854
rect 520706 305778 521262 306334
rect 524426 309498 524982 310054
rect 523130 294938 523366 295174
rect 523130 294618 523366 294854
rect 520706 269778 521262 270334
rect 524426 273498 524982 274054
rect 523130 258938 523366 259174
rect 523130 258618 523366 258854
rect 520706 233778 521262 234334
rect 524426 237498 524982 238054
rect 523130 222938 523366 223174
rect 523130 222618 523366 222854
rect 520706 197778 521262 198334
rect 524426 201498 524982 202054
rect 523130 186938 523366 187174
rect 523130 186618 523366 186854
rect 520706 161778 521262 162334
rect 524426 165498 524982 166054
rect 523130 150938 523366 151174
rect 523130 150618 523366 150854
rect 520706 125778 521262 126334
rect 524426 129498 524982 130054
rect 523130 114938 523366 115174
rect 523130 114618 523366 114854
rect 520706 89778 521262 90334
rect 524426 93498 524982 94054
rect 523130 78938 523366 79174
rect 523130 78618 523366 78854
rect 520706 53778 521262 54334
rect 524426 57498 524982 58054
rect 523130 42938 523366 43174
rect 523130 42618 523366 42854
rect 520706 17778 521262 18334
rect 524426 21498 524982 22054
rect 523130 6938 523366 7174
rect 523130 6618 523366 6854
rect 520706 -4742 521262 -4186
rect 524426 -5702 524982 -5146
rect 528146 710042 528702 710598
rect 528146 673218 528702 673774
rect 528146 637218 528702 637774
rect 528146 601218 528702 601774
rect 528146 565218 528702 565774
rect 528146 529218 528702 529774
rect 528146 493218 528702 493774
rect 528146 457218 528702 457774
rect 528146 421218 528702 421774
rect 528146 385218 528702 385774
rect 528146 349218 528702 349774
rect 528146 313218 528702 313774
rect 528146 277218 528702 277774
rect 528146 241218 528702 241774
rect 528146 205218 528702 205774
rect 528146 169218 528702 169774
rect 528146 133218 528702 133774
rect 528146 97218 528702 97774
rect 528146 61218 528702 61774
rect 528146 25218 528702 25774
rect 528146 -6662 528702 -6106
rect 531866 711002 532422 711558
rect 531866 676938 532422 677494
rect 531866 640938 532422 641494
rect 531866 604938 532422 605494
rect 531866 568938 532422 569494
rect 531866 532938 532422 533494
rect 531866 496938 532422 497494
rect 531866 460938 532422 461494
rect 531866 424938 532422 425494
rect 531866 388938 532422 389494
rect 531866 352938 532422 353494
rect 541826 704282 542382 704838
rect 541826 686898 542382 687454
rect 541826 650898 542382 651454
rect 541826 614898 542382 615454
rect 541826 578898 542382 579454
rect 541826 542898 542382 543454
rect 541826 506898 542382 507454
rect 541826 470898 542382 471454
rect 541826 434898 542382 435454
rect 541826 398898 542382 399454
rect 541826 362898 542382 363454
rect 538490 327218 538726 327454
rect 538490 326898 538726 327134
rect 541826 326898 542382 327454
rect 531866 316938 532422 317494
rect 538490 291218 538726 291454
rect 538490 290898 538726 291134
rect 541826 290898 542382 291454
rect 531866 280938 532422 281494
rect 538490 255218 538726 255454
rect 538490 254898 538726 255134
rect 541826 254898 542382 255454
rect 531866 244938 532422 245494
rect 538490 219218 538726 219454
rect 538490 218898 538726 219134
rect 541826 218898 542382 219454
rect 531866 208938 532422 209494
rect 538490 183218 538726 183454
rect 538490 182898 538726 183134
rect 541826 182898 542382 183454
rect 531866 172938 532422 173494
rect 538490 147218 538726 147454
rect 538490 146898 538726 147134
rect 541826 146898 542382 147454
rect 531866 136938 532422 137494
rect 538490 111218 538726 111454
rect 538490 110898 538726 111134
rect 541826 110898 542382 111454
rect 531866 100938 532422 101494
rect 538490 75218 538726 75454
rect 538490 74898 538726 75134
rect 541826 74898 542382 75454
rect 531866 64938 532422 65494
rect 538490 39218 538726 39454
rect 538490 38898 538726 39134
rect 541826 38898 542382 39454
rect 531866 28938 532422 29494
rect 531866 -7622 532422 -7066
rect 541826 2898 542382 3454
rect 541826 -902 542382 -346
rect 545546 705242 546102 705798
rect 545546 690618 546102 691174
rect 545546 654618 546102 655174
rect 545546 618618 546102 619174
rect 545546 582618 546102 583174
rect 545546 546618 546102 547174
rect 545546 510618 546102 511174
rect 545546 474618 546102 475174
rect 545546 438618 546102 439174
rect 545546 402618 546102 403174
rect 545546 366618 546102 367174
rect 545546 330618 546102 331174
rect 545546 294618 546102 295174
rect 545546 258618 546102 259174
rect 545546 222618 546102 223174
rect 545546 186618 546102 187174
rect 545546 150618 546102 151174
rect 545546 114618 546102 115174
rect 545546 78618 546102 79174
rect 545546 42618 546102 43174
rect 545546 6618 546102 7174
rect 545546 -1862 546102 -1306
rect 549266 706202 549822 706758
rect 549266 694338 549822 694894
rect 549266 658338 549822 658894
rect 549266 622338 549822 622894
rect 549266 586338 549822 586894
rect 549266 550338 549822 550894
rect 549266 514338 549822 514894
rect 549266 478338 549822 478894
rect 549266 442338 549822 442894
rect 549266 406338 549822 406894
rect 549266 370338 549822 370894
rect 549266 334338 549822 334894
rect 549266 298338 549822 298894
rect 549266 262338 549822 262894
rect 549266 226338 549822 226894
rect 549266 190338 549822 190894
rect 549266 154338 549822 154894
rect 549266 118338 549822 118894
rect 549266 82338 549822 82894
rect 549266 46338 549822 46894
rect 549266 10338 549822 10894
rect 549266 -2822 549822 -2266
rect 552986 707162 553542 707718
rect 552986 698058 553542 698614
rect 552986 662058 553542 662614
rect 552986 626058 553542 626614
rect 552986 590058 553542 590614
rect 552986 554058 553542 554614
rect 552986 518058 553542 518614
rect 552986 482058 553542 482614
rect 552986 446058 553542 446614
rect 552986 410058 553542 410614
rect 552986 374058 553542 374614
rect 552986 338058 553542 338614
rect 556706 708122 557262 708678
rect 556706 665778 557262 666334
rect 556706 629778 557262 630334
rect 556706 593778 557262 594334
rect 556706 557778 557262 558334
rect 556706 521778 557262 522334
rect 556706 485778 557262 486334
rect 556706 449778 557262 450334
rect 556706 413778 557262 414334
rect 556706 377778 557262 378334
rect 556706 341778 557262 342334
rect 553850 330938 554086 331174
rect 553850 330618 554086 330854
rect 552986 302058 553542 302614
rect 556706 305778 557262 306334
rect 553850 294938 554086 295174
rect 553850 294618 554086 294854
rect 552986 266058 553542 266614
rect 556706 269778 557262 270334
rect 553850 258938 554086 259174
rect 553850 258618 554086 258854
rect 552986 230058 553542 230614
rect 556706 233778 557262 234334
rect 553850 222938 554086 223174
rect 553850 222618 554086 222854
rect 552986 194058 553542 194614
rect 556706 197778 557262 198334
rect 553850 186938 554086 187174
rect 553850 186618 554086 186854
rect 552986 158058 553542 158614
rect 556706 161778 557262 162334
rect 553850 150938 554086 151174
rect 553850 150618 554086 150854
rect 552986 122058 553542 122614
rect 556706 125778 557262 126334
rect 553850 114938 554086 115174
rect 553850 114618 554086 114854
rect 552986 86058 553542 86614
rect 556706 89778 557262 90334
rect 553850 78938 554086 79174
rect 553850 78618 554086 78854
rect 552986 50058 553542 50614
rect 556706 53778 557262 54334
rect 553850 42938 554086 43174
rect 553850 42618 554086 42854
rect 552986 14058 553542 14614
rect 556706 17778 557262 18334
rect 553850 6938 554086 7174
rect 553850 6618 554086 6854
rect 552986 -3782 553542 -3226
rect 556706 -4742 557262 -4186
rect 560426 709082 560982 709638
rect 560426 669498 560982 670054
rect 560426 633498 560982 634054
rect 560426 597498 560982 598054
rect 560426 561498 560982 562054
rect 560426 525498 560982 526054
rect 560426 489498 560982 490054
rect 560426 453498 560982 454054
rect 560426 417498 560982 418054
rect 560426 381498 560982 382054
rect 560426 345498 560982 346054
rect 560426 309498 560982 310054
rect 560426 273498 560982 274054
rect 560426 237498 560982 238054
rect 560426 201498 560982 202054
rect 560426 165498 560982 166054
rect 560426 129498 560982 130054
rect 560426 93498 560982 94054
rect 560426 57498 560982 58054
rect 560426 21498 560982 22054
rect 560426 -5702 560982 -5146
rect 564146 710042 564702 710598
rect 564146 673218 564702 673774
rect 564146 637218 564702 637774
rect 564146 601218 564702 601774
rect 564146 565218 564702 565774
rect 564146 529218 564702 529774
rect 564146 493218 564702 493774
rect 564146 457218 564702 457774
rect 564146 421218 564702 421774
rect 564146 385218 564702 385774
rect 564146 349218 564702 349774
rect 564146 313218 564702 313774
rect 564146 277218 564702 277774
rect 564146 241218 564702 241774
rect 564146 205218 564702 205774
rect 564146 169218 564702 169774
rect 564146 133218 564702 133774
rect 564146 97218 564702 97774
rect 564146 61218 564702 61774
rect 564146 25218 564702 25774
rect 564146 -6662 564702 -6106
rect 567866 711002 568422 711558
rect 567866 676938 568422 677494
rect 567866 640938 568422 641494
rect 567866 604938 568422 605494
rect 567866 568938 568422 569494
rect 567866 532938 568422 533494
rect 567866 496938 568422 497494
rect 567866 460938 568422 461494
rect 567866 424938 568422 425494
rect 567866 388938 568422 389494
rect 567866 352938 568422 353494
rect 577826 704282 578382 704838
rect 577826 686898 578382 687454
rect 577826 650898 578382 651454
rect 577826 614898 578382 615454
rect 577826 578898 578382 579454
rect 577826 542898 578382 543454
rect 577826 506898 578382 507454
rect 577826 470898 578382 471454
rect 577826 434898 578382 435454
rect 577826 398898 578382 399454
rect 577826 362898 578382 363454
rect 569210 327218 569446 327454
rect 569210 326898 569446 327134
rect 577826 326898 578382 327454
rect 567866 316938 568422 317494
rect 569210 291218 569446 291454
rect 569210 290898 569446 291134
rect 577826 290898 578382 291454
rect 567866 280938 568422 281494
rect 569210 255218 569446 255454
rect 569210 254898 569446 255134
rect 577826 254898 578382 255454
rect 567866 244938 568422 245494
rect 569210 219218 569446 219454
rect 569210 218898 569446 219134
rect 577826 218898 578382 219454
rect 567866 208938 568422 209494
rect 569210 183218 569446 183454
rect 569210 182898 569446 183134
rect 577826 182898 578382 183454
rect 567866 172938 568422 173494
rect 569210 147218 569446 147454
rect 569210 146898 569446 147134
rect 577826 146898 578382 147454
rect 567866 136938 568422 137494
rect 569210 111218 569446 111454
rect 569210 110898 569446 111134
rect 577826 110898 578382 111454
rect 567866 100938 568422 101494
rect 569210 75218 569446 75454
rect 569210 74898 569446 75134
rect 577826 74898 578382 75454
rect 567866 64938 568422 65494
rect 569210 39218 569446 39454
rect 569210 38898 569446 39134
rect 577826 38898 578382 39454
rect 567866 28938 568422 29494
rect 567866 -7622 568422 -7066
rect 577826 2898 578382 3454
rect 577826 -902 578382 -346
rect 592062 711002 592618 711558
rect 591102 710042 591658 710598
rect 590142 709082 590698 709638
rect 589182 708122 589738 708678
rect 588222 707162 588778 707718
rect 587262 706202 587818 706758
rect 581546 705242 582102 705798
rect 586302 705242 586858 705798
rect 581546 690618 582102 691174
rect 581546 654618 582102 655174
rect 581546 618618 582102 619174
rect 581546 582618 582102 583174
rect 581546 546618 582102 547174
rect 581546 510618 582102 511174
rect 581546 474618 582102 475174
rect 581546 438618 582102 439174
rect 581546 402618 582102 403174
rect 581546 366618 582102 367174
rect 581546 330618 582102 331174
rect 581546 294618 582102 295174
rect 581546 258618 582102 259174
rect 581546 222618 582102 223174
rect 581546 186618 582102 187174
rect 581546 150618 582102 151174
rect 581546 114618 582102 115174
rect 581546 78618 582102 79174
rect 581546 42618 582102 43174
rect 581546 6618 582102 7174
rect 585342 704282 585898 704838
rect 585342 686898 585898 687454
rect 585342 650898 585898 651454
rect 585342 614898 585898 615454
rect 585342 578898 585898 579454
rect 585342 542898 585898 543454
rect 585342 506898 585898 507454
rect 585342 470898 585898 471454
rect 585342 434898 585898 435454
rect 585342 398898 585898 399454
rect 585342 362898 585898 363454
rect 585342 326898 585898 327454
rect 585342 290898 585898 291454
rect 585342 254898 585898 255454
rect 585342 218898 585898 219454
rect 585342 182898 585898 183454
rect 585342 146898 585898 147454
rect 585342 110898 585898 111454
rect 585342 74898 585898 75454
rect 585342 38898 585898 39454
rect 585342 2898 585898 3454
rect 585342 -902 585898 -346
rect 586302 690618 586858 691174
rect 586302 654618 586858 655174
rect 586302 618618 586858 619174
rect 586302 582618 586858 583174
rect 586302 546618 586858 547174
rect 586302 510618 586858 511174
rect 586302 474618 586858 475174
rect 586302 438618 586858 439174
rect 586302 402618 586858 403174
rect 586302 366618 586858 367174
rect 586302 330618 586858 331174
rect 586302 294618 586858 295174
rect 586302 258618 586858 259174
rect 586302 222618 586858 223174
rect 586302 186618 586858 187174
rect 586302 150618 586858 151174
rect 586302 114618 586858 115174
rect 586302 78618 586858 79174
rect 586302 42618 586858 43174
rect 586302 6618 586858 7174
rect 581546 -1862 582102 -1306
rect 586302 -1862 586858 -1306
rect 587262 694338 587818 694894
rect 587262 658338 587818 658894
rect 587262 622338 587818 622894
rect 587262 586338 587818 586894
rect 587262 550338 587818 550894
rect 587262 514338 587818 514894
rect 587262 478338 587818 478894
rect 587262 442338 587818 442894
rect 587262 406338 587818 406894
rect 587262 370338 587818 370894
rect 587262 334338 587818 334894
rect 587262 298338 587818 298894
rect 587262 262338 587818 262894
rect 587262 226338 587818 226894
rect 587262 190338 587818 190894
rect 587262 154338 587818 154894
rect 587262 118338 587818 118894
rect 587262 82338 587818 82894
rect 587262 46338 587818 46894
rect 587262 10338 587818 10894
rect 587262 -2822 587818 -2266
rect 588222 698058 588778 698614
rect 588222 662058 588778 662614
rect 588222 626058 588778 626614
rect 588222 590058 588778 590614
rect 588222 554058 588778 554614
rect 588222 518058 588778 518614
rect 588222 482058 588778 482614
rect 588222 446058 588778 446614
rect 588222 410058 588778 410614
rect 588222 374058 588778 374614
rect 588222 338058 588778 338614
rect 588222 302058 588778 302614
rect 588222 266058 588778 266614
rect 588222 230058 588778 230614
rect 588222 194058 588778 194614
rect 588222 158058 588778 158614
rect 588222 122058 588778 122614
rect 588222 86058 588778 86614
rect 588222 50058 588778 50614
rect 588222 14058 588778 14614
rect 588222 -3782 588778 -3226
rect 589182 665778 589738 666334
rect 589182 629778 589738 630334
rect 589182 593778 589738 594334
rect 589182 557778 589738 558334
rect 589182 521778 589738 522334
rect 589182 485778 589738 486334
rect 589182 449778 589738 450334
rect 589182 413778 589738 414334
rect 589182 377778 589738 378334
rect 589182 341778 589738 342334
rect 589182 305778 589738 306334
rect 589182 269778 589738 270334
rect 589182 233778 589738 234334
rect 589182 197778 589738 198334
rect 589182 161778 589738 162334
rect 589182 125778 589738 126334
rect 589182 89778 589738 90334
rect 589182 53778 589738 54334
rect 589182 17778 589738 18334
rect 589182 -4742 589738 -4186
rect 590142 669498 590698 670054
rect 590142 633498 590698 634054
rect 590142 597498 590698 598054
rect 590142 561498 590698 562054
rect 590142 525498 590698 526054
rect 590142 489498 590698 490054
rect 590142 453498 590698 454054
rect 590142 417498 590698 418054
rect 590142 381498 590698 382054
rect 590142 345498 590698 346054
rect 590142 309498 590698 310054
rect 590142 273498 590698 274054
rect 590142 237498 590698 238054
rect 590142 201498 590698 202054
rect 590142 165498 590698 166054
rect 590142 129498 590698 130054
rect 590142 93498 590698 94054
rect 590142 57498 590698 58054
rect 590142 21498 590698 22054
rect 590142 -5702 590698 -5146
rect 591102 673218 591658 673774
rect 591102 637218 591658 637774
rect 591102 601218 591658 601774
rect 591102 565218 591658 565774
rect 591102 529218 591658 529774
rect 591102 493218 591658 493774
rect 591102 457218 591658 457774
rect 591102 421218 591658 421774
rect 591102 385218 591658 385774
rect 591102 349218 591658 349774
rect 591102 313218 591658 313774
rect 591102 277218 591658 277774
rect 591102 241218 591658 241774
rect 591102 205218 591658 205774
rect 591102 169218 591658 169774
rect 591102 133218 591658 133774
rect 591102 97218 591658 97774
rect 591102 61218 591658 61774
rect 591102 25218 591658 25774
rect 591102 -6662 591658 -6106
rect 592062 676938 592618 677494
rect 592062 640938 592618 641494
rect 592062 604938 592618 605494
rect 592062 568938 592618 569494
rect 592062 532938 592618 533494
rect 592062 496938 592618 497494
rect 592062 460938 592618 461494
rect 592062 424938 592618 425494
rect 592062 388938 592618 389494
rect 592062 352938 592618 353494
rect 592062 316938 592618 317494
rect 592062 280938 592618 281494
rect 592062 244938 592618 245494
rect 592062 208938 592618 209494
rect 592062 172938 592618 173494
rect 592062 136938 592618 137494
rect 592062 100938 592618 101494
rect 592062 64938 592618 65494
rect 592062 28938 592618 29494
rect 592062 -7622 592618 -7066
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711002 -8694 711558
rect -8138 711002 27866 711558
rect 28422 711002 63866 711558
rect 64422 711002 99866 711558
rect 100422 711002 135866 711558
rect 136422 711002 171866 711558
rect 172422 711002 207866 711558
rect 208422 711002 243866 711558
rect 244422 711002 279866 711558
rect 280422 711002 315866 711558
rect 316422 711002 351866 711558
rect 352422 711002 387866 711558
rect 388422 711002 423866 711558
rect 424422 711002 459866 711558
rect 460422 711002 495866 711558
rect 496422 711002 531866 711558
rect 532422 711002 567866 711558
rect 568422 711002 592062 711558
rect 592618 711002 592650 711558
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710042 -7734 710598
rect -7178 710042 24146 710598
rect 24702 710042 60146 710598
rect 60702 710042 96146 710598
rect 96702 710042 132146 710598
rect 132702 710042 168146 710598
rect 168702 710042 204146 710598
rect 204702 710042 240146 710598
rect 240702 710042 276146 710598
rect 276702 710042 312146 710598
rect 312702 710042 348146 710598
rect 348702 710042 384146 710598
rect 384702 710042 420146 710598
rect 420702 710042 456146 710598
rect 456702 710042 492146 710598
rect 492702 710042 528146 710598
rect 528702 710042 564146 710598
rect 564702 710042 591102 710598
rect 591658 710042 591690 710598
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709082 -6774 709638
rect -6218 709082 20426 709638
rect 20982 709082 56426 709638
rect 56982 709082 92426 709638
rect 92982 709082 128426 709638
rect 128982 709082 164426 709638
rect 164982 709082 200426 709638
rect 200982 709082 236426 709638
rect 236982 709082 272426 709638
rect 272982 709082 308426 709638
rect 308982 709082 344426 709638
rect 344982 709082 380426 709638
rect 380982 709082 416426 709638
rect 416982 709082 452426 709638
rect 452982 709082 488426 709638
rect 488982 709082 524426 709638
rect 524982 709082 560426 709638
rect 560982 709082 590142 709638
rect 590698 709082 590730 709638
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708122 -5814 708678
rect -5258 708122 16706 708678
rect 17262 708122 52706 708678
rect 53262 708122 88706 708678
rect 89262 708122 124706 708678
rect 125262 708122 160706 708678
rect 161262 708122 196706 708678
rect 197262 708122 232706 708678
rect 233262 708122 268706 708678
rect 269262 708122 304706 708678
rect 305262 708122 340706 708678
rect 341262 708122 376706 708678
rect 377262 708122 412706 708678
rect 413262 708122 448706 708678
rect 449262 708122 484706 708678
rect 485262 708122 520706 708678
rect 521262 708122 556706 708678
rect 557262 708122 589182 708678
rect 589738 708122 589770 708678
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707162 -4854 707718
rect -4298 707162 12986 707718
rect 13542 707162 48986 707718
rect 49542 707162 84986 707718
rect 85542 707162 120986 707718
rect 121542 707162 156986 707718
rect 157542 707162 192986 707718
rect 193542 707162 228986 707718
rect 229542 707162 264986 707718
rect 265542 707162 300986 707718
rect 301542 707162 336986 707718
rect 337542 707162 372986 707718
rect 373542 707162 408986 707718
rect 409542 707162 444986 707718
rect 445542 707162 480986 707718
rect 481542 707162 516986 707718
rect 517542 707162 552986 707718
rect 553542 707162 588222 707718
rect 588778 707162 588810 707718
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706202 -3894 706758
rect -3338 706202 9266 706758
rect 9822 706202 45266 706758
rect 45822 706202 81266 706758
rect 81822 706202 117266 706758
rect 117822 706202 153266 706758
rect 153822 706202 189266 706758
rect 189822 706202 225266 706758
rect 225822 706202 261266 706758
rect 261822 706202 297266 706758
rect 297822 706202 333266 706758
rect 333822 706202 369266 706758
rect 369822 706202 405266 706758
rect 405822 706202 441266 706758
rect 441822 706202 477266 706758
rect 477822 706202 513266 706758
rect 513822 706202 549266 706758
rect 549822 706202 587262 706758
rect 587818 706202 587850 706758
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705242 -2934 705798
rect -2378 705242 5546 705798
rect 6102 705242 41546 705798
rect 42102 705242 77546 705798
rect 78102 705242 113546 705798
rect 114102 705242 149546 705798
rect 150102 705242 185546 705798
rect 186102 705242 221546 705798
rect 222102 705242 257546 705798
rect 258102 705242 293546 705798
rect 294102 705242 329546 705798
rect 330102 705242 365546 705798
rect 366102 705242 401546 705798
rect 402102 705242 437546 705798
rect 438102 705242 473546 705798
rect 474102 705242 509546 705798
rect 510102 705242 545546 705798
rect 546102 705242 581546 705798
rect 582102 705242 586302 705798
rect 586858 705242 586890 705798
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704282 -1974 704838
rect -1418 704282 1826 704838
rect 2382 704282 37826 704838
rect 38382 704282 73826 704838
rect 74382 704282 109826 704838
rect 110382 704282 145826 704838
rect 146382 704282 181826 704838
rect 182382 704282 217826 704838
rect 218382 704282 253826 704838
rect 254382 704282 289826 704838
rect 290382 704282 325826 704838
rect 326382 704282 361826 704838
rect 362382 704282 397826 704838
rect 398382 704282 433826 704838
rect 434382 704282 469826 704838
rect 470382 704282 505826 704838
rect 506382 704282 541826 704838
rect 542382 704282 577826 704838
rect 578382 704282 585342 704838
rect 585898 704282 585930 704838
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698058 -4854 698614
rect -4298 698058 12986 698614
rect 13542 698058 48986 698614
rect 49542 698058 84986 698614
rect 85542 698058 120986 698614
rect 121542 698058 156986 698614
rect 157542 698058 192986 698614
rect 193542 698058 228986 698614
rect 229542 698058 264986 698614
rect 265542 698058 300986 698614
rect 301542 698058 336986 698614
rect 337542 698058 372986 698614
rect 373542 698058 408986 698614
rect 409542 698058 444986 698614
rect 445542 698058 480986 698614
rect 481542 698058 516986 698614
rect 517542 698058 552986 698614
rect 553542 698058 588222 698614
rect 588778 698058 592650 698614
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694338 -3894 694894
rect -3338 694338 9266 694894
rect 9822 694338 45266 694894
rect 45822 694338 81266 694894
rect 81822 694338 117266 694894
rect 117822 694338 153266 694894
rect 153822 694338 189266 694894
rect 189822 694338 225266 694894
rect 225822 694338 261266 694894
rect 261822 694338 297266 694894
rect 297822 694338 333266 694894
rect 333822 694338 369266 694894
rect 369822 694338 405266 694894
rect 405822 694338 441266 694894
rect 441822 694338 477266 694894
rect 477822 694338 513266 694894
rect 513822 694338 549266 694894
rect 549822 694338 587262 694894
rect 587818 694338 592650 694894
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690618 -2934 691174
rect -2378 690618 5546 691174
rect 6102 690618 41546 691174
rect 42102 690618 77546 691174
rect 78102 690618 113546 691174
rect 114102 690618 149546 691174
rect 150102 690618 185546 691174
rect 186102 690618 221546 691174
rect 222102 690618 257546 691174
rect 258102 690618 293546 691174
rect 294102 690618 329546 691174
rect 330102 690618 365546 691174
rect 366102 690618 401546 691174
rect 402102 690618 437546 691174
rect 438102 690618 473546 691174
rect 474102 690618 509546 691174
rect 510102 690618 545546 691174
rect 546102 690618 581546 691174
rect 582102 690618 586302 691174
rect 586858 690618 592650 691174
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 686898 -1974 687454
rect -1418 686898 1826 687454
rect 2382 686898 37826 687454
rect 38382 686898 73826 687454
rect 74382 686898 109826 687454
rect 110382 686898 145826 687454
rect 146382 686898 181826 687454
rect 182382 686898 217826 687454
rect 218382 686898 253826 687454
rect 254382 686898 289826 687454
rect 290382 686898 325826 687454
rect 326382 686898 361826 687454
rect 362382 686898 397826 687454
rect 398382 686898 433826 687454
rect 434382 686898 469826 687454
rect 470382 686898 505826 687454
rect 506382 686898 541826 687454
rect 542382 686898 577826 687454
rect 578382 686898 585342 687454
rect 585898 686898 592650 687454
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 676938 -8694 677494
rect -8138 676938 27866 677494
rect 28422 676938 63866 677494
rect 64422 676938 99866 677494
rect 100422 676938 135866 677494
rect 136422 676938 171866 677494
rect 172422 676938 207866 677494
rect 208422 676938 243866 677494
rect 244422 676938 279866 677494
rect 280422 676938 315866 677494
rect 316422 676938 351866 677494
rect 352422 676938 387866 677494
rect 388422 676938 423866 677494
rect 424422 676938 459866 677494
rect 460422 676938 495866 677494
rect 496422 676938 531866 677494
rect 532422 676938 567866 677494
rect 568422 676938 592062 677494
rect 592618 676938 592650 677494
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673218 -7734 673774
rect -7178 673218 24146 673774
rect 24702 673218 60146 673774
rect 60702 673218 96146 673774
rect 96702 673218 132146 673774
rect 132702 673218 168146 673774
rect 168702 673218 204146 673774
rect 204702 673218 240146 673774
rect 240702 673218 276146 673774
rect 276702 673218 312146 673774
rect 312702 673218 348146 673774
rect 348702 673218 384146 673774
rect 384702 673218 420146 673774
rect 420702 673218 456146 673774
rect 456702 673218 492146 673774
rect 492702 673218 528146 673774
rect 528702 673218 564146 673774
rect 564702 673218 591102 673774
rect 591658 673218 592650 673774
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669498 -6774 670054
rect -6218 669498 20426 670054
rect 20982 669498 56426 670054
rect 56982 669498 92426 670054
rect 92982 669498 128426 670054
rect 128982 669498 164426 670054
rect 164982 669498 200426 670054
rect 200982 669498 236426 670054
rect 236982 669498 272426 670054
rect 272982 669498 308426 670054
rect 308982 669498 344426 670054
rect 344982 669498 380426 670054
rect 380982 669498 416426 670054
rect 416982 669498 452426 670054
rect 452982 669498 488426 670054
rect 488982 669498 524426 670054
rect 524982 669498 560426 670054
rect 560982 669498 590142 670054
rect 590698 669498 592650 670054
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 665778 -5814 666334
rect -5258 665778 16706 666334
rect 17262 665778 52706 666334
rect 53262 665778 88706 666334
rect 89262 665778 124706 666334
rect 125262 665778 160706 666334
rect 161262 665778 196706 666334
rect 197262 665778 232706 666334
rect 233262 665778 268706 666334
rect 269262 665778 304706 666334
rect 305262 665778 340706 666334
rect 341262 665778 376706 666334
rect 377262 665778 412706 666334
rect 413262 665778 448706 666334
rect 449262 665778 484706 666334
rect 485262 665778 520706 666334
rect 521262 665778 556706 666334
rect 557262 665778 589182 666334
rect 589738 665778 592650 666334
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662058 -4854 662614
rect -4298 662058 12986 662614
rect 13542 662058 48986 662614
rect 49542 662058 84986 662614
rect 85542 662058 120986 662614
rect 121542 662058 156986 662614
rect 157542 662058 192986 662614
rect 193542 662058 228986 662614
rect 229542 662058 264986 662614
rect 265542 662058 300986 662614
rect 301542 662058 336986 662614
rect 337542 662058 372986 662614
rect 373542 662058 408986 662614
rect 409542 662058 444986 662614
rect 445542 662058 480986 662614
rect 481542 662058 516986 662614
rect 517542 662058 552986 662614
rect 553542 662058 588222 662614
rect 588778 662058 592650 662614
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658338 -3894 658894
rect -3338 658338 9266 658894
rect 9822 658338 45266 658894
rect 45822 658338 81266 658894
rect 81822 658338 117266 658894
rect 117822 658338 153266 658894
rect 153822 658338 189266 658894
rect 189822 658338 225266 658894
rect 225822 658338 261266 658894
rect 261822 658338 297266 658894
rect 297822 658338 333266 658894
rect 333822 658338 369266 658894
rect 369822 658338 405266 658894
rect 405822 658338 441266 658894
rect 441822 658338 477266 658894
rect 477822 658338 513266 658894
rect 513822 658338 549266 658894
rect 549822 658338 587262 658894
rect 587818 658338 592650 658894
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654618 -2934 655174
rect -2378 654618 5546 655174
rect 6102 654618 41546 655174
rect 42102 654618 77546 655174
rect 78102 654618 113546 655174
rect 114102 654618 149546 655174
rect 150102 654618 185546 655174
rect 186102 654618 221546 655174
rect 222102 654618 257546 655174
rect 258102 654618 293546 655174
rect 294102 654618 329546 655174
rect 330102 654618 365546 655174
rect 366102 654618 401546 655174
rect 402102 654618 437546 655174
rect 438102 654618 473546 655174
rect 474102 654618 509546 655174
rect 510102 654618 545546 655174
rect 546102 654618 581546 655174
rect 582102 654618 586302 655174
rect 586858 654618 592650 655174
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 650898 -1974 651454
rect -1418 650898 1826 651454
rect 2382 650898 37826 651454
rect 38382 650898 73826 651454
rect 74382 650898 109826 651454
rect 110382 650898 145826 651454
rect 146382 650898 181826 651454
rect 182382 650898 217826 651454
rect 218382 650898 253826 651454
rect 254382 650898 289826 651454
rect 290382 650898 325826 651454
rect 326382 650898 361826 651454
rect 362382 650898 397826 651454
rect 398382 650898 433826 651454
rect 434382 650898 469826 651454
rect 470382 650898 505826 651454
rect 506382 650898 541826 651454
rect 542382 650898 577826 651454
rect 578382 650898 585342 651454
rect 585898 650898 592650 651454
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 640938 -8694 641494
rect -8138 640938 27866 641494
rect 28422 640938 63866 641494
rect 64422 640938 99866 641494
rect 100422 640938 135866 641494
rect 136422 640938 171866 641494
rect 172422 640938 207866 641494
rect 208422 640938 243866 641494
rect 244422 640938 279866 641494
rect 280422 640938 315866 641494
rect 316422 640938 351866 641494
rect 352422 640938 387866 641494
rect 388422 640938 423866 641494
rect 424422 640938 459866 641494
rect 460422 640938 495866 641494
rect 496422 640938 531866 641494
rect 532422 640938 567866 641494
rect 568422 640938 592062 641494
rect 592618 640938 592650 641494
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637218 -7734 637774
rect -7178 637218 24146 637774
rect 24702 637218 60146 637774
rect 60702 637218 96146 637774
rect 96702 637218 132146 637774
rect 132702 637218 168146 637774
rect 168702 637218 204146 637774
rect 204702 637218 240146 637774
rect 240702 637218 276146 637774
rect 276702 637218 312146 637774
rect 312702 637218 348146 637774
rect 348702 637218 384146 637774
rect 384702 637218 420146 637774
rect 420702 637218 456146 637774
rect 456702 637218 492146 637774
rect 492702 637218 528146 637774
rect 528702 637218 564146 637774
rect 564702 637218 591102 637774
rect 591658 637218 592650 637774
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633498 -6774 634054
rect -6218 633498 20426 634054
rect 20982 633498 56426 634054
rect 56982 633498 92426 634054
rect 92982 633498 128426 634054
rect 128982 633498 164426 634054
rect 164982 633498 200426 634054
rect 200982 633498 236426 634054
rect 236982 633498 272426 634054
rect 272982 633498 308426 634054
rect 308982 633498 344426 634054
rect 344982 633498 380426 634054
rect 380982 633498 416426 634054
rect 416982 633498 452426 634054
rect 452982 633498 488426 634054
rect 488982 633498 524426 634054
rect 524982 633498 560426 634054
rect 560982 633498 590142 634054
rect 590698 633498 592650 634054
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 629778 -5814 630334
rect -5258 629778 16706 630334
rect 17262 629778 52706 630334
rect 53262 629778 88706 630334
rect 89262 629778 124706 630334
rect 125262 629778 160706 630334
rect 161262 629778 196706 630334
rect 197262 629778 232706 630334
rect 233262 629778 268706 630334
rect 269262 629778 304706 630334
rect 305262 629778 340706 630334
rect 341262 629778 376706 630334
rect 377262 629778 412706 630334
rect 413262 629778 448706 630334
rect 449262 629778 484706 630334
rect 485262 629778 520706 630334
rect 521262 629778 556706 630334
rect 557262 629778 589182 630334
rect 589738 629778 592650 630334
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626058 -4854 626614
rect -4298 626058 12986 626614
rect 13542 626058 48986 626614
rect 49542 626058 84986 626614
rect 85542 626058 120986 626614
rect 121542 626058 156986 626614
rect 157542 626058 192986 626614
rect 193542 626058 228986 626614
rect 229542 626058 264986 626614
rect 265542 626058 300986 626614
rect 301542 626058 336986 626614
rect 337542 626058 372986 626614
rect 373542 626058 408986 626614
rect 409542 626058 444986 626614
rect 445542 626058 480986 626614
rect 481542 626058 516986 626614
rect 517542 626058 552986 626614
rect 553542 626058 588222 626614
rect 588778 626058 592650 626614
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622338 -3894 622894
rect -3338 622338 9266 622894
rect 9822 622338 45266 622894
rect 45822 622338 81266 622894
rect 81822 622338 117266 622894
rect 117822 622338 153266 622894
rect 153822 622338 189266 622894
rect 189822 622338 225266 622894
rect 225822 622338 261266 622894
rect 261822 622338 297266 622894
rect 297822 622338 333266 622894
rect 333822 622338 369266 622894
rect 369822 622338 405266 622894
rect 405822 622338 441266 622894
rect 441822 622338 477266 622894
rect 477822 622338 513266 622894
rect 513822 622338 549266 622894
rect 549822 622338 587262 622894
rect 587818 622338 592650 622894
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618618 -2934 619174
rect -2378 618618 5546 619174
rect 6102 618618 41546 619174
rect 42102 618618 77546 619174
rect 78102 618618 113546 619174
rect 114102 618618 149546 619174
rect 150102 618618 185546 619174
rect 186102 618618 221546 619174
rect 222102 618618 257546 619174
rect 258102 618618 293546 619174
rect 294102 618618 329546 619174
rect 330102 618618 365546 619174
rect 366102 618618 401546 619174
rect 402102 618618 437546 619174
rect 438102 618618 473546 619174
rect 474102 618618 509546 619174
rect 510102 618618 545546 619174
rect 546102 618618 581546 619174
rect 582102 618618 586302 619174
rect 586858 618618 592650 619174
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 614898 -1974 615454
rect -1418 614898 1826 615454
rect 2382 614898 37826 615454
rect 38382 614898 73826 615454
rect 74382 614898 109826 615454
rect 110382 614898 145826 615454
rect 146382 614898 181826 615454
rect 182382 614898 217826 615454
rect 218382 614898 253826 615454
rect 254382 614898 289826 615454
rect 290382 614898 325826 615454
rect 326382 614898 361826 615454
rect 362382 614898 397826 615454
rect 398382 614898 433826 615454
rect 434382 614898 469826 615454
rect 470382 614898 505826 615454
rect 506382 614898 541826 615454
rect 542382 614898 577826 615454
rect 578382 614898 585342 615454
rect 585898 614898 592650 615454
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 604938 -8694 605494
rect -8138 604938 27866 605494
rect 28422 604938 63866 605494
rect 64422 604938 99866 605494
rect 100422 604938 135866 605494
rect 136422 604938 171866 605494
rect 172422 604938 207866 605494
rect 208422 604938 243866 605494
rect 244422 604938 279866 605494
rect 280422 604938 315866 605494
rect 316422 604938 351866 605494
rect 352422 604938 387866 605494
rect 388422 604938 423866 605494
rect 424422 604938 459866 605494
rect 460422 604938 495866 605494
rect 496422 604938 531866 605494
rect 532422 604938 567866 605494
rect 568422 604938 592062 605494
rect 592618 604938 592650 605494
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601218 -7734 601774
rect -7178 601218 24146 601774
rect 24702 601218 60146 601774
rect 60702 601218 96146 601774
rect 96702 601218 132146 601774
rect 132702 601218 168146 601774
rect 168702 601218 204146 601774
rect 204702 601218 240146 601774
rect 240702 601218 276146 601774
rect 276702 601218 312146 601774
rect 312702 601218 348146 601774
rect 348702 601218 384146 601774
rect 384702 601218 420146 601774
rect 420702 601218 456146 601774
rect 456702 601218 492146 601774
rect 492702 601218 528146 601774
rect 528702 601218 564146 601774
rect 564702 601218 591102 601774
rect 591658 601218 592650 601774
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597498 -6774 598054
rect -6218 597498 20426 598054
rect 20982 597498 56426 598054
rect 56982 597498 92426 598054
rect 92982 597498 128426 598054
rect 128982 597498 164426 598054
rect 164982 597498 200426 598054
rect 200982 597498 236426 598054
rect 236982 597498 272426 598054
rect 272982 597498 308426 598054
rect 308982 597498 344426 598054
rect 344982 597498 380426 598054
rect 380982 597498 416426 598054
rect 416982 597498 452426 598054
rect 452982 597498 488426 598054
rect 488982 597498 524426 598054
rect 524982 597498 560426 598054
rect 560982 597498 590142 598054
rect 590698 597498 592650 598054
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 593778 -5814 594334
rect -5258 593778 16706 594334
rect 17262 593778 52706 594334
rect 53262 593778 88706 594334
rect 89262 593778 124706 594334
rect 125262 593778 160706 594334
rect 161262 593778 196706 594334
rect 197262 593778 232706 594334
rect 233262 593778 268706 594334
rect 269262 593778 304706 594334
rect 305262 593778 340706 594334
rect 341262 593778 376706 594334
rect 377262 593778 412706 594334
rect 413262 593778 448706 594334
rect 449262 593778 484706 594334
rect 485262 593778 520706 594334
rect 521262 593778 556706 594334
rect 557262 593778 589182 594334
rect 589738 593778 592650 594334
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590058 -4854 590614
rect -4298 590058 12986 590614
rect 13542 590058 48986 590614
rect 49542 590058 84986 590614
rect 85542 590058 120986 590614
rect 121542 590058 156986 590614
rect 157542 590058 192986 590614
rect 193542 590058 228986 590614
rect 229542 590058 264986 590614
rect 265542 590058 300986 590614
rect 301542 590058 336986 590614
rect 337542 590058 372986 590614
rect 373542 590058 408986 590614
rect 409542 590058 444986 590614
rect 445542 590058 480986 590614
rect 481542 590058 516986 590614
rect 517542 590058 552986 590614
rect 553542 590058 588222 590614
rect 588778 590058 592650 590614
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586338 -3894 586894
rect -3338 586338 9266 586894
rect 9822 586338 45266 586894
rect 45822 586338 81266 586894
rect 81822 586338 117266 586894
rect 117822 586338 153266 586894
rect 153822 586338 189266 586894
rect 189822 586338 225266 586894
rect 225822 586338 261266 586894
rect 261822 586338 297266 586894
rect 297822 586338 333266 586894
rect 333822 586338 369266 586894
rect 369822 586338 405266 586894
rect 405822 586338 441266 586894
rect 441822 586338 477266 586894
rect 477822 586338 513266 586894
rect 513822 586338 549266 586894
rect 549822 586338 587262 586894
rect 587818 586338 592650 586894
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582618 -2934 583174
rect -2378 582618 5546 583174
rect 6102 582618 41546 583174
rect 42102 582618 77546 583174
rect 78102 582618 113546 583174
rect 114102 582618 149546 583174
rect 150102 582618 185546 583174
rect 186102 582618 221546 583174
rect 222102 582618 257546 583174
rect 258102 582618 293546 583174
rect 294102 582618 329546 583174
rect 330102 582618 365546 583174
rect 366102 582618 401546 583174
rect 402102 582618 437546 583174
rect 438102 582618 473546 583174
rect 474102 582618 509546 583174
rect 510102 582618 545546 583174
rect 546102 582618 581546 583174
rect 582102 582618 586302 583174
rect 586858 582618 592650 583174
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 578898 -1974 579454
rect -1418 578898 1826 579454
rect 2382 578898 37826 579454
rect 38382 578898 73826 579454
rect 74382 578898 109826 579454
rect 110382 578898 145826 579454
rect 146382 578898 181826 579454
rect 182382 578898 217826 579454
rect 218382 578898 253826 579454
rect 254382 578898 289826 579454
rect 290382 578898 325826 579454
rect 326382 578898 361826 579454
rect 362382 578898 397826 579454
rect 398382 578898 433826 579454
rect 434382 578898 469826 579454
rect 470382 578898 505826 579454
rect 506382 578898 541826 579454
rect 542382 578898 577826 579454
rect 578382 578898 585342 579454
rect 585898 578898 592650 579454
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 568938 -8694 569494
rect -8138 568938 27866 569494
rect 28422 568938 63866 569494
rect 64422 568938 99866 569494
rect 100422 568938 135866 569494
rect 136422 568938 171866 569494
rect 172422 568938 207866 569494
rect 208422 568938 243866 569494
rect 244422 568938 279866 569494
rect 280422 568938 315866 569494
rect 316422 568938 351866 569494
rect 352422 568938 387866 569494
rect 388422 568938 423866 569494
rect 424422 568938 459866 569494
rect 460422 568938 495866 569494
rect 496422 568938 531866 569494
rect 532422 568938 567866 569494
rect 568422 568938 592062 569494
rect 592618 568938 592650 569494
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565218 -7734 565774
rect -7178 565218 24146 565774
rect 24702 565218 60146 565774
rect 60702 565218 96146 565774
rect 96702 565218 132146 565774
rect 132702 565218 168146 565774
rect 168702 565218 204146 565774
rect 204702 565218 240146 565774
rect 240702 565218 276146 565774
rect 276702 565218 312146 565774
rect 312702 565218 348146 565774
rect 348702 565218 384146 565774
rect 384702 565218 420146 565774
rect 420702 565218 456146 565774
rect 456702 565218 492146 565774
rect 492702 565218 528146 565774
rect 528702 565218 564146 565774
rect 564702 565218 591102 565774
rect 591658 565218 592650 565774
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561498 -6774 562054
rect -6218 561498 20426 562054
rect 20982 561498 56426 562054
rect 56982 561498 92426 562054
rect 92982 561498 128426 562054
rect 128982 561498 164426 562054
rect 164982 561498 200426 562054
rect 200982 561498 236426 562054
rect 236982 561498 272426 562054
rect 272982 561498 308426 562054
rect 308982 561498 344426 562054
rect 344982 561498 380426 562054
rect 380982 561498 416426 562054
rect 416982 561498 452426 562054
rect 452982 561498 488426 562054
rect 488982 561498 524426 562054
rect 524982 561498 560426 562054
rect 560982 561498 590142 562054
rect 590698 561498 592650 562054
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 557778 -5814 558334
rect -5258 557778 16706 558334
rect 17262 557778 52706 558334
rect 53262 557778 88706 558334
rect 89262 557778 124706 558334
rect 125262 557778 160706 558334
rect 161262 557778 196706 558334
rect 197262 557778 232706 558334
rect 233262 557778 268706 558334
rect 269262 557778 304706 558334
rect 305262 557778 340706 558334
rect 341262 557778 376706 558334
rect 377262 557778 412706 558334
rect 413262 557778 448706 558334
rect 449262 557778 484706 558334
rect 485262 557778 520706 558334
rect 521262 557778 556706 558334
rect 557262 557778 589182 558334
rect 589738 557778 592650 558334
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554058 -4854 554614
rect -4298 554058 12986 554614
rect 13542 554058 48986 554614
rect 49542 554058 84986 554614
rect 85542 554058 120986 554614
rect 121542 554058 156986 554614
rect 157542 554058 192986 554614
rect 193542 554058 228986 554614
rect 229542 554058 264986 554614
rect 265542 554058 300986 554614
rect 301542 554058 336986 554614
rect 337542 554058 372986 554614
rect 373542 554058 408986 554614
rect 409542 554058 444986 554614
rect 445542 554058 480986 554614
rect 481542 554058 516986 554614
rect 517542 554058 552986 554614
rect 553542 554058 588222 554614
rect 588778 554058 592650 554614
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550338 -3894 550894
rect -3338 550338 9266 550894
rect 9822 550338 45266 550894
rect 45822 550338 81266 550894
rect 81822 550338 117266 550894
rect 117822 550338 153266 550894
rect 153822 550338 189266 550894
rect 189822 550338 225266 550894
rect 225822 550338 261266 550894
rect 261822 550338 297266 550894
rect 297822 550338 333266 550894
rect 333822 550338 369266 550894
rect 369822 550338 405266 550894
rect 405822 550338 441266 550894
rect 441822 550338 477266 550894
rect 477822 550338 513266 550894
rect 513822 550338 549266 550894
rect 549822 550338 587262 550894
rect 587818 550338 592650 550894
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546618 -2934 547174
rect -2378 546618 5546 547174
rect 6102 546618 41546 547174
rect 42102 546618 77546 547174
rect 78102 546618 113546 547174
rect 114102 546618 149546 547174
rect 150102 546618 185546 547174
rect 186102 546618 221546 547174
rect 222102 546618 257546 547174
rect 258102 546618 293546 547174
rect 294102 546618 329546 547174
rect 330102 546618 365546 547174
rect 366102 546618 401546 547174
rect 402102 546618 437546 547174
rect 438102 546618 473546 547174
rect 474102 546618 509546 547174
rect 510102 546618 545546 547174
rect 546102 546618 581546 547174
rect 582102 546618 586302 547174
rect 586858 546618 592650 547174
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 542898 -1974 543454
rect -1418 542898 1826 543454
rect 2382 542898 37826 543454
rect 38382 542898 73826 543454
rect 74382 542898 109826 543454
rect 110382 542898 145826 543454
rect 146382 542898 181826 543454
rect 182382 542898 217826 543454
rect 218382 542898 253826 543454
rect 254382 542898 289826 543454
rect 290382 542898 325826 543454
rect 326382 542898 361826 543454
rect 362382 542898 397826 543454
rect 398382 542898 433826 543454
rect 434382 542898 469826 543454
rect 470382 542898 505826 543454
rect 506382 542898 541826 543454
rect 542382 542898 577826 543454
rect 578382 542898 585342 543454
rect 585898 542898 592650 543454
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 532938 -8694 533494
rect -8138 532938 27866 533494
rect 28422 532938 63866 533494
rect 64422 532938 99866 533494
rect 100422 532938 135866 533494
rect 136422 532938 171866 533494
rect 172422 532938 207866 533494
rect 208422 532938 243866 533494
rect 244422 532938 279866 533494
rect 280422 532938 315866 533494
rect 316422 532938 351866 533494
rect 352422 532938 387866 533494
rect 388422 532938 423866 533494
rect 424422 532938 459866 533494
rect 460422 532938 495866 533494
rect 496422 532938 531866 533494
rect 532422 532938 567866 533494
rect 568422 532938 592062 533494
rect 592618 532938 592650 533494
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529218 -7734 529774
rect -7178 529218 24146 529774
rect 24702 529218 60146 529774
rect 60702 529218 96146 529774
rect 96702 529218 132146 529774
rect 132702 529218 168146 529774
rect 168702 529218 204146 529774
rect 204702 529218 240146 529774
rect 240702 529218 276146 529774
rect 276702 529218 312146 529774
rect 312702 529218 348146 529774
rect 348702 529218 384146 529774
rect 384702 529218 420146 529774
rect 420702 529218 456146 529774
rect 456702 529218 492146 529774
rect 492702 529218 528146 529774
rect 528702 529218 564146 529774
rect 564702 529218 591102 529774
rect 591658 529218 592650 529774
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525498 -6774 526054
rect -6218 525498 20426 526054
rect 20982 525498 56426 526054
rect 56982 525498 92426 526054
rect 92982 525498 128426 526054
rect 128982 525498 164426 526054
rect 164982 525498 200426 526054
rect 200982 525498 236426 526054
rect 236982 525498 272426 526054
rect 272982 525498 308426 526054
rect 308982 525498 344426 526054
rect 344982 525498 380426 526054
rect 380982 525498 416426 526054
rect 416982 525498 452426 526054
rect 452982 525498 488426 526054
rect 488982 525498 524426 526054
rect 524982 525498 560426 526054
rect 560982 525498 590142 526054
rect 590698 525498 592650 526054
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 521778 -5814 522334
rect -5258 521778 16706 522334
rect 17262 521778 52706 522334
rect 53262 521778 88706 522334
rect 89262 521778 124706 522334
rect 125262 521778 160706 522334
rect 161262 521778 196706 522334
rect 197262 521778 232706 522334
rect 233262 521778 268706 522334
rect 269262 521778 304706 522334
rect 305262 521778 340706 522334
rect 341262 521778 376706 522334
rect 377262 521778 412706 522334
rect 413262 521778 448706 522334
rect 449262 521778 484706 522334
rect 485262 521778 520706 522334
rect 521262 521778 556706 522334
rect 557262 521778 589182 522334
rect 589738 521778 592650 522334
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518058 -4854 518614
rect -4298 518058 12986 518614
rect 13542 518058 48986 518614
rect 49542 518058 84986 518614
rect 85542 518058 120986 518614
rect 121542 518058 156986 518614
rect 157542 518058 192986 518614
rect 193542 518058 228986 518614
rect 229542 518058 264986 518614
rect 265542 518058 300986 518614
rect 301542 518058 336986 518614
rect 337542 518058 372986 518614
rect 373542 518058 408986 518614
rect 409542 518058 444986 518614
rect 445542 518058 480986 518614
rect 481542 518058 516986 518614
rect 517542 518058 552986 518614
rect 553542 518058 588222 518614
rect 588778 518058 592650 518614
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514338 -3894 514894
rect -3338 514338 9266 514894
rect 9822 514338 45266 514894
rect 45822 514338 81266 514894
rect 81822 514338 117266 514894
rect 117822 514338 153266 514894
rect 153822 514338 189266 514894
rect 189822 514338 225266 514894
rect 225822 514338 261266 514894
rect 261822 514338 297266 514894
rect 297822 514338 333266 514894
rect 333822 514338 369266 514894
rect 369822 514338 405266 514894
rect 405822 514338 441266 514894
rect 441822 514338 477266 514894
rect 477822 514338 513266 514894
rect 513822 514338 549266 514894
rect 549822 514338 587262 514894
rect 587818 514338 592650 514894
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510618 -2934 511174
rect -2378 510618 5546 511174
rect 6102 510618 41546 511174
rect 42102 510618 77546 511174
rect 78102 510618 113546 511174
rect 114102 510618 149546 511174
rect 150102 510618 185546 511174
rect 186102 510618 221546 511174
rect 222102 510618 257546 511174
rect 258102 510618 293546 511174
rect 294102 510618 329546 511174
rect 330102 510618 365546 511174
rect 366102 510618 401546 511174
rect 402102 510618 437546 511174
rect 438102 510618 473546 511174
rect 474102 510618 509546 511174
rect 510102 510618 545546 511174
rect 546102 510618 581546 511174
rect 582102 510618 586302 511174
rect 586858 510618 592650 511174
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 506898 -1974 507454
rect -1418 506898 1826 507454
rect 2382 506898 37826 507454
rect 38382 506898 73826 507454
rect 74382 506898 109826 507454
rect 110382 506898 145826 507454
rect 146382 506898 181826 507454
rect 182382 506898 217826 507454
rect 218382 506898 253826 507454
rect 254382 506898 289826 507454
rect 290382 506898 325826 507454
rect 326382 506898 361826 507454
rect 362382 506898 397826 507454
rect 398382 506898 433826 507454
rect 434382 506898 469826 507454
rect 470382 506898 505826 507454
rect 506382 506898 541826 507454
rect 542382 506898 577826 507454
rect 578382 506898 585342 507454
rect 585898 506898 592650 507454
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 496938 -8694 497494
rect -8138 496938 27866 497494
rect 28422 496938 63866 497494
rect 64422 496938 99866 497494
rect 100422 496938 135866 497494
rect 136422 496938 171866 497494
rect 172422 496938 207866 497494
rect 208422 496938 243866 497494
rect 244422 496938 279866 497494
rect 280422 496938 315866 497494
rect 316422 496938 351866 497494
rect 352422 496938 387866 497494
rect 388422 496938 423866 497494
rect 424422 496938 459866 497494
rect 460422 496938 495866 497494
rect 496422 496938 531866 497494
rect 532422 496938 567866 497494
rect 568422 496938 592062 497494
rect 592618 496938 592650 497494
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493218 -7734 493774
rect -7178 493218 24146 493774
rect 24702 493218 60146 493774
rect 60702 493218 96146 493774
rect 96702 493218 132146 493774
rect 132702 493218 168146 493774
rect 168702 493218 204146 493774
rect 204702 493218 240146 493774
rect 240702 493218 276146 493774
rect 276702 493218 312146 493774
rect 312702 493218 348146 493774
rect 348702 493218 384146 493774
rect 384702 493218 420146 493774
rect 420702 493218 456146 493774
rect 456702 493218 492146 493774
rect 492702 493218 528146 493774
rect 528702 493218 564146 493774
rect 564702 493218 591102 493774
rect 591658 493218 592650 493774
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489498 -6774 490054
rect -6218 489498 20426 490054
rect 20982 489498 56426 490054
rect 56982 489498 92426 490054
rect 92982 489498 128426 490054
rect 128982 489498 164426 490054
rect 164982 489498 200426 490054
rect 200982 489498 236426 490054
rect 236982 489498 272426 490054
rect 272982 489498 308426 490054
rect 308982 489498 344426 490054
rect 344982 489498 380426 490054
rect 380982 489498 416426 490054
rect 416982 489498 452426 490054
rect 452982 489498 488426 490054
rect 488982 489498 524426 490054
rect 524982 489498 560426 490054
rect 560982 489498 590142 490054
rect 590698 489498 592650 490054
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 485778 -5814 486334
rect -5258 485778 16706 486334
rect 17262 485778 52706 486334
rect 53262 485778 88706 486334
rect 89262 485778 124706 486334
rect 125262 485778 160706 486334
rect 161262 485778 196706 486334
rect 197262 485778 232706 486334
rect 233262 485778 268706 486334
rect 269262 485778 304706 486334
rect 305262 485778 340706 486334
rect 341262 485778 376706 486334
rect 377262 485778 412706 486334
rect 413262 485778 448706 486334
rect 449262 485778 484706 486334
rect 485262 485778 520706 486334
rect 521262 485778 556706 486334
rect 557262 485778 589182 486334
rect 589738 485778 592650 486334
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482058 -4854 482614
rect -4298 482058 12986 482614
rect 13542 482058 48986 482614
rect 49542 482058 84986 482614
rect 85542 482058 120986 482614
rect 121542 482058 156986 482614
rect 157542 482058 192986 482614
rect 193542 482058 228986 482614
rect 229542 482058 264986 482614
rect 265542 482058 300986 482614
rect 301542 482058 336986 482614
rect 337542 482058 372986 482614
rect 373542 482058 408986 482614
rect 409542 482058 444986 482614
rect 445542 482058 480986 482614
rect 481542 482058 516986 482614
rect 517542 482058 552986 482614
rect 553542 482058 588222 482614
rect 588778 482058 592650 482614
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478338 -3894 478894
rect -3338 478338 9266 478894
rect 9822 478338 45266 478894
rect 45822 478338 81266 478894
rect 81822 478338 117266 478894
rect 117822 478338 153266 478894
rect 153822 478338 189266 478894
rect 189822 478338 225266 478894
rect 225822 478338 261266 478894
rect 261822 478338 297266 478894
rect 297822 478338 333266 478894
rect 333822 478338 369266 478894
rect 369822 478338 405266 478894
rect 405822 478338 441266 478894
rect 441822 478338 477266 478894
rect 477822 478338 513266 478894
rect 513822 478338 549266 478894
rect 549822 478338 587262 478894
rect 587818 478338 592650 478894
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474618 -2934 475174
rect -2378 474618 5546 475174
rect 6102 474618 41546 475174
rect 42102 474618 77546 475174
rect 78102 474618 113546 475174
rect 114102 474618 149546 475174
rect 150102 474618 185546 475174
rect 186102 474618 221546 475174
rect 222102 474618 257546 475174
rect 258102 474618 293546 475174
rect 294102 474618 329546 475174
rect 330102 474618 365546 475174
rect 366102 474618 401546 475174
rect 402102 474618 437546 475174
rect 438102 474618 473546 475174
rect 474102 474618 509546 475174
rect 510102 474618 545546 475174
rect 546102 474618 581546 475174
rect 582102 474618 586302 475174
rect 586858 474618 592650 475174
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 470898 -1974 471454
rect -1418 470898 1826 471454
rect 2382 470898 37826 471454
rect 38382 470898 73826 471454
rect 74382 470898 109826 471454
rect 110382 470898 145826 471454
rect 146382 470898 181826 471454
rect 182382 470898 217826 471454
rect 218382 470898 253826 471454
rect 254382 470898 289826 471454
rect 290382 470898 325826 471454
rect 326382 470898 361826 471454
rect 362382 470898 397826 471454
rect 398382 470898 433826 471454
rect 434382 470898 469826 471454
rect 470382 470898 505826 471454
rect 506382 470898 541826 471454
rect 542382 470898 577826 471454
rect 578382 470898 585342 471454
rect 585898 470898 592650 471454
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 460938 -8694 461494
rect -8138 460938 27866 461494
rect 28422 460938 63866 461494
rect 64422 460938 99866 461494
rect 100422 460938 135866 461494
rect 136422 460938 171866 461494
rect 172422 460938 207866 461494
rect 208422 460938 243866 461494
rect 244422 460938 279866 461494
rect 280422 460938 315866 461494
rect 316422 460938 351866 461494
rect 352422 460938 387866 461494
rect 388422 460938 423866 461494
rect 424422 460938 459866 461494
rect 460422 460938 495866 461494
rect 496422 460938 531866 461494
rect 532422 460938 567866 461494
rect 568422 460938 592062 461494
rect 592618 460938 592650 461494
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457218 -7734 457774
rect -7178 457218 24146 457774
rect 24702 457218 60146 457774
rect 60702 457218 96146 457774
rect 96702 457218 132146 457774
rect 132702 457218 168146 457774
rect 168702 457218 204146 457774
rect 204702 457218 240146 457774
rect 240702 457218 276146 457774
rect 276702 457218 312146 457774
rect 312702 457218 348146 457774
rect 348702 457218 384146 457774
rect 384702 457218 420146 457774
rect 420702 457218 456146 457774
rect 456702 457218 492146 457774
rect 492702 457218 528146 457774
rect 528702 457218 564146 457774
rect 564702 457218 591102 457774
rect 591658 457218 592650 457774
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453498 -6774 454054
rect -6218 453498 20426 454054
rect 20982 453498 56426 454054
rect 56982 453498 92426 454054
rect 92982 453498 128426 454054
rect 128982 453498 164426 454054
rect 164982 453498 200426 454054
rect 200982 453498 236426 454054
rect 236982 453498 272426 454054
rect 272982 453498 308426 454054
rect 308982 453498 344426 454054
rect 344982 453498 380426 454054
rect 380982 453498 416426 454054
rect 416982 453498 452426 454054
rect 452982 453498 488426 454054
rect 488982 453498 524426 454054
rect 524982 453498 560426 454054
rect 560982 453498 590142 454054
rect 590698 453498 592650 454054
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 449778 -5814 450334
rect -5258 449778 16706 450334
rect 17262 449778 52706 450334
rect 53262 449778 88706 450334
rect 89262 449778 124706 450334
rect 125262 449778 160706 450334
rect 161262 449778 196706 450334
rect 197262 449778 232706 450334
rect 233262 449778 268706 450334
rect 269262 449778 304706 450334
rect 305262 449778 340706 450334
rect 341262 449778 376706 450334
rect 377262 449778 412706 450334
rect 413262 449778 448706 450334
rect 449262 449778 484706 450334
rect 485262 449778 520706 450334
rect 521262 449778 556706 450334
rect 557262 449778 589182 450334
rect 589738 449778 592650 450334
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446058 -4854 446614
rect -4298 446058 12986 446614
rect 13542 446058 48986 446614
rect 49542 446058 84986 446614
rect 85542 446058 120986 446614
rect 121542 446058 156986 446614
rect 157542 446058 192986 446614
rect 193542 446058 228986 446614
rect 229542 446058 264986 446614
rect 265542 446058 300986 446614
rect 301542 446058 336986 446614
rect 337542 446058 372986 446614
rect 373542 446058 408986 446614
rect 409542 446058 444986 446614
rect 445542 446058 480986 446614
rect 481542 446058 516986 446614
rect 517542 446058 552986 446614
rect 553542 446058 588222 446614
rect 588778 446058 592650 446614
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442338 -3894 442894
rect -3338 442338 9266 442894
rect 9822 442338 45266 442894
rect 45822 442338 81266 442894
rect 81822 442338 117266 442894
rect 117822 442338 153266 442894
rect 153822 442338 189266 442894
rect 189822 442338 225266 442894
rect 225822 442338 261266 442894
rect 261822 442338 297266 442894
rect 297822 442338 333266 442894
rect 333822 442338 369266 442894
rect 369822 442338 405266 442894
rect 405822 442338 441266 442894
rect 441822 442338 477266 442894
rect 477822 442338 513266 442894
rect 513822 442338 549266 442894
rect 549822 442338 587262 442894
rect 587818 442338 592650 442894
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438618 -2934 439174
rect -2378 438618 5546 439174
rect 6102 438618 41546 439174
rect 42102 438618 77546 439174
rect 78102 438618 113546 439174
rect 114102 438618 149546 439174
rect 150102 438618 185546 439174
rect 186102 438618 221546 439174
rect 222102 438618 257546 439174
rect 258102 438618 293546 439174
rect 294102 438618 329546 439174
rect 330102 438618 365546 439174
rect 366102 438618 401546 439174
rect 402102 438618 437546 439174
rect 438102 438618 473546 439174
rect 474102 438618 509546 439174
rect 510102 438618 545546 439174
rect 546102 438618 581546 439174
rect 582102 438618 586302 439174
rect 586858 438618 592650 439174
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 434898 -1974 435454
rect -1418 434898 1826 435454
rect 2382 434898 37826 435454
rect 38382 434898 73826 435454
rect 74382 434898 109826 435454
rect 110382 434898 145826 435454
rect 146382 434898 181826 435454
rect 182382 434898 217826 435454
rect 218382 434898 253826 435454
rect 254382 434898 289826 435454
rect 290382 434898 325826 435454
rect 326382 434898 361826 435454
rect 362382 434898 397826 435454
rect 398382 434898 433826 435454
rect 434382 434898 469826 435454
rect 470382 434898 505826 435454
rect 506382 434898 541826 435454
rect 542382 434898 577826 435454
rect 578382 434898 585342 435454
rect 585898 434898 592650 435454
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 424938 -8694 425494
rect -8138 424938 27866 425494
rect 28422 424938 63866 425494
rect 64422 424938 99866 425494
rect 100422 424938 135866 425494
rect 136422 424938 171866 425494
rect 172422 424938 207866 425494
rect 208422 424938 243866 425494
rect 244422 424938 279866 425494
rect 280422 424938 315866 425494
rect 316422 424938 351866 425494
rect 352422 424938 387866 425494
rect 388422 424938 423866 425494
rect 424422 424938 459866 425494
rect 460422 424938 495866 425494
rect 496422 424938 531866 425494
rect 532422 424938 567866 425494
rect 568422 424938 592062 425494
rect 592618 424938 592650 425494
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421218 -7734 421774
rect -7178 421218 24146 421774
rect 24702 421218 60146 421774
rect 60702 421218 96146 421774
rect 96702 421218 132146 421774
rect 132702 421218 168146 421774
rect 168702 421218 204146 421774
rect 204702 421218 240146 421774
rect 240702 421218 276146 421774
rect 276702 421218 312146 421774
rect 312702 421218 348146 421774
rect 348702 421218 384146 421774
rect 384702 421218 420146 421774
rect 420702 421218 456146 421774
rect 456702 421218 492146 421774
rect 492702 421218 528146 421774
rect 528702 421218 564146 421774
rect 564702 421218 591102 421774
rect 591658 421218 592650 421774
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417498 -6774 418054
rect -6218 417498 20426 418054
rect 20982 417498 56426 418054
rect 56982 417498 92426 418054
rect 92982 417498 128426 418054
rect 128982 417498 164426 418054
rect 164982 417498 200426 418054
rect 200982 417498 236426 418054
rect 236982 417498 272426 418054
rect 272982 417498 308426 418054
rect 308982 417498 344426 418054
rect 344982 417498 380426 418054
rect 380982 417498 416426 418054
rect 416982 417498 452426 418054
rect 452982 417498 488426 418054
rect 488982 417498 524426 418054
rect 524982 417498 560426 418054
rect 560982 417498 590142 418054
rect 590698 417498 592650 418054
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 413778 -5814 414334
rect -5258 413778 16706 414334
rect 17262 413778 52706 414334
rect 53262 413778 88706 414334
rect 89262 413778 124706 414334
rect 125262 413778 160706 414334
rect 161262 413778 196706 414334
rect 197262 413778 232706 414334
rect 233262 413778 268706 414334
rect 269262 413778 304706 414334
rect 305262 413778 340706 414334
rect 341262 413778 376706 414334
rect 377262 413778 412706 414334
rect 413262 413778 448706 414334
rect 449262 413778 484706 414334
rect 485262 413778 520706 414334
rect 521262 413778 556706 414334
rect 557262 413778 589182 414334
rect 589738 413778 592650 414334
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410058 -4854 410614
rect -4298 410058 12986 410614
rect 13542 410058 48986 410614
rect 49542 410058 84986 410614
rect 85542 410058 120986 410614
rect 121542 410058 156986 410614
rect 157542 410058 192986 410614
rect 193542 410058 228986 410614
rect 229542 410058 264986 410614
rect 265542 410058 300986 410614
rect 301542 410058 336986 410614
rect 337542 410058 372986 410614
rect 373542 410058 408986 410614
rect 409542 410058 444986 410614
rect 445542 410058 480986 410614
rect 481542 410058 516986 410614
rect 517542 410058 552986 410614
rect 553542 410058 588222 410614
rect 588778 410058 592650 410614
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406338 -3894 406894
rect -3338 406338 9266 406894
rect 9822 406338 45266 406894
rect 45822 406338 81266 406894
rect 81822 406338 117266 406894
rect 117822 406338 153266 406894
rect 153822 406338 189266 406894
rect 189822 406338 225266 406894
rect 225822 406338 261266 406894
rect 261822 406338 297266 406894
rect 297822 406338 333266 406894
rect 333822 406338 369266 406894
rect 369822 406338 405266 406894
rect 405822 406338 441266 406894
rect 441822 406338 477266 406894
rect 477822 406338 513266 406894
rect 513822 406338 549266 406894
rect 549822 406338 587262 406894
rect 587818 406338 592650 406894
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402618 -2934 403174
rect -2378 402618 5546 403174
rect 6102 402618 41546 403174
rect 42102 402618 77546 403174
rect 78102 402618 113546 403174
rect 114102 402618 149546 403174
rect 150102 402618 185546 403174
rect 186102 402618 221546 403174
rect 222102 402618 257546 403174
rect 258102 402618 293546 403174
rect 294102 402618 329546 403174
rect 330102 402618 365546 403174
rect 366102 402618 401546 403174
rect 402102 402618 437546 403174
rect 438102 402618 473546 403174
rect 474102 402618 509546 403174
rect 510102 402618 545546 403174
rect 546102 402618 581546 403174
rect 582102 402618 586302 403174
rect 586858 402618 592650 403174
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 398898 -1974 399454
rect -1418 398898 1826 399454
rect 2382 398898 37826 399454
rect 38382 398898 73826 399454
rect 74382 398898 109826 399454
rect 110382 398898 145826 399454
rect 146382 398898 181826 399454
rect 182382 398898 217826 399454
rect 218382 398898 253826 399454
rect 254382 398898 289826 399454
rect 290382 398898 325826 399454
rect 326382 398898 361826 399454
rect 362382 398898 397826 399454
rect 398382 398898 433826 399454
rect 434382 398898 469826 399454
rect 470382 398898 505826 399454
rect 506382 398898 541826 399454
rect 542382 398898 577826 399454
rect 578382 398898 585342 399454
rect 585898 398898 592650 399454
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 388938 -8694 389494
rect -8138 388938 27866 389494
rect 28422 388938 63866 389494
rect 64422 388938 99866 389494
rect 100422 388938 135866 389494
rect 136422 388938 171866 389494
rect 172422 388938 207866 389494
rect 208422 388938 243866 389494
rect 244422 388938 279866 389494
rect 280422 388938 315866 389494
rect 316422 388938 351866 389494
rect 352422 388938 387866 389494
rect 388422 388938 423866 389494
rect 424422 388938 459866 389494
rect 460422 388938 495866 389494
rect 496422 388938 531866 389494
rect 532422 388938 567866 389494
rect 568422 388938 592062 389494
rect 592618 388938 592650 389494
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385218 -7734 385774
rect -7178 385218 24146 385774
rect 24702 385218 60146 385774
rect 60702 385218 96146 385774
rect 96702 385218 132146 385774
rect 132702 385218 168146 385774
rect 168702 385218 204146 385774
rect 204702 385218 240146 385774
rect 240702 385218 276146 385774
rect 276702 385218 312146 385774
rect 312702 385218 348146 385774
rect 348702 385218 384146 385774
rect 384702 385218 420146 385774
rect 420702 385218 456146 385774
rect 456702 385218 492146 385774
rect 492702 385218 528146 385774
rect 528702 385218 564146 385774
rect 564702 385218 591102 385774
rect 591658 385218 592650 385774
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381498 -6774 382054
rect -6218 381498 20426 382054
rect 20982 381498 56426 382054
rect 56982 381498 92426 382054
rect 92982 381498 128426 382054
rect 128982 381498 164426 382054
rect 164982 381498 200426 382054
rect 200982 381498 236426 382054
rect 236982 381498 272426 382054
rect 272982 381498 308426 382054
rect 308982 381498 344426 382054
rect 344982 381498 380426 382054
rect 380982 381498 416426 382054
rect 416982 381498 452426 382054
rect 452982 381498 488426 382054
rect 488982 381498 524426 382054
rect 524982 381498 560426 382054
rect 560982 381498 590142 382054
rect 590698 381498 592650 382054
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 377778 -5814 378334
rect -5258 377778 16706 378334
rect 17262 377778 52706 378334
rect 53262 377778 88706 378334
rect 89262 377778 124706 378334
rect 125262 377778 160706 378334
rect 161262 377778 196706 378334
rect 197262 377778 232706 378334
rect 233262 377778 268706 378334
rect 269262 377778 304706 378334
rect 305262 377778 340706 378334
rect 341262 377778 376706 378334
rect 377262 377778 412706 378334
rect 413262 377778 448706 378334
rect 449262 377778 484706 378334
rect 485262 377778 520706 378334
rect 521262 377778 556706 378334
rect 557262 377778 589182 378334
rect 589738 377778 592650 378334
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374058 -4854 374614
rect -4298 374058 12986 374614
rect 13542 374058 48986 374614
rect 49542 374058 84986 374614
rect 85542 374058 120986 374614
rect 121542 374058 156986 374614
rect 157542 374058 192986 374614
rect 193542 374058 228986 374614
rect 229542 374058 264986 374614
rect 265542 374058 300986 374614
rect 301542 374058 336986 374614
rect 337542 374058 372986 374614
rect 373542 374058 408986 374614
rect 409542 374058 444986 374614
rect 445542 374058 480986 374614
rect 481542 374058 516986 374614
rect 517542 374058 552986 374614
rect 553542 374058 588222 374614
rect 588778 374058 592650 374614
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370338 -3894 370894
rect -3338 370338 9266 370894
rect 9822 370338 45266 370894
rect 45822 370338 81266 370894
rect 81822 370338 117266 370894
rect 117822 370338 153266 370894
rect 153822 370338 189266 370894
rect 189822 370338 225266 370894
rect 225822 370338 261266 370894
rect 261822 370338 297266 370894
rect 297822 370338 333266 370894
rect 333822 370338 369266 370894
rect 369822 370338 405266 370894
rect 405822 370338 441266 370894
rect 441822 370338 477266 370894
rect 477822 370338 513266 370894
rect 513822 370338 549266 370894
rect 549822 370338 587262 370894
rect 587818 370338 592650 370894
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366618 -2934 367174
rect -2378 366618 5546 367174
rect 6102 366618 41546 367174
rect 42102 366618 77546 367174
rect 78102 366618 113546 367174
rect 114102 366618 149546 367174
rect 150102 366618 185546 367174
rect 186102 366618 221546 367174
rect 222102 366618 257546 367174
rect 258102 366618 293546 367174
rect 294102 366618 329546 367174
rect 330102 366618 365546 367174
rect 366102 366618 401546 367174
rect 402102 366618 437546 367174
rect 438102 366618 473546 367174
rect 474102 366618 509546 367174
rect 510102 366618 545546 367174
rect 546102 366618 581546 367174
rect 582102 366618 586302 367174
rect 586858 366618 592650 367174
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 362898 -1974 363454
rect -1418 362898 1826 363454
rect 2382 362898 37826 363454
rect 38382 362898 73826 363454
rect 74382 362898 109826 363454
rect 110382 362898 145826 363454
rect 146382 362898 181826 363454
rect 182382 362898 217826 363454
rect 218382 362898 253826 363454
rect 254382 362898 289826 363454
rect 290382 362898 325826 363454
rect 326382 362898 361826 363454
rect 362382 362898 397826 363454
rect 398382 362898 433826 363454
rect 434382 362898 469826 363454
rect 470382 362898 505826 363454
rect 506382 362898 541826 363454
rect 542382 362898 577826 363454
rect 578382 362898 585342 363454
rect 585898 362898 592650 363454
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 352938 -8694 353494
rect -8138 352938 27866 353494
rect 28422 352938 63866 353494
rect 64422 352938 99866 353494
rect 100422 352938 135866 353494
rect 136422 352938 171866 353494
rect 172422 352938 207866 353494
rect 208422 352938 243866 353494
rect 244422 352938 279866 353494
rect 280422 352938 315866 353494
rect 316422 352938 351866 353494
rect 352422 352938 387866 353494
rect 388422 352938 423866 353494
rect 424422 352938 459866 353494
rect 460422 352938 495866 353494
rect 496422 352938 531866 353494
rect 532422 352938 567866 353494
rect 568422 352938 592062 353494
rect 592618 352938 592650 353494
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349218 -7734 349774
rect -7178 349218 24146 349774
rect 24702 349218 60146 349774
rect 60702 349218 96146 349774
rect 96702 349218 132146 349774
rect 132702 349218 168146 349774
rect 168702 349218 204146 349774
rect 204702 349218 240146 349774
rect 240702 349218 276146 349774
rect 276702 349218 312146 349774
rect 312702 349218 348146 349774
rect 348702 349218 384146 349774
rect 384702 349218 420146 349774
rect 420702 349218 456146 349774
rect 456702 349218 528146 349774
rect 528702 349218 564146 349774
rect 564702 349218 591102 349774
rect 591658 349218 592650 349774
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345498 -6774 346054
rect -6218 345498 20426 346054
rect 20982 345498 56426 346054
rect 56982 345498 128426 346054
rect 128982 345498 164426 346054
rect 164982 345498 236426 346054
rect 236982 345498 272426 346054
rect 272982 345498 344426 346054
rect 344982 345498 380426 346054
rect 380982 345498 416426 346054
rect 416982 345498 452426 346054
rect 452982 345498 488426 346054
rect 488982 345498 524426 346054
rect 524982 345498 560426 346054
rect 560982 345498 590142 346054
rect 590698 345498 592650 346054
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 341778 -5814 342334
rect -5258 341778 16706 342334
rect 17262 341778 52706 342334
rect 53262 341778 88706 342334
rect 89262 341778 124706 342334
rect 125262 341778 160706 342334
rect 161262 341778 196706 342334
rect 197262 341778 232706 342334
rect 233262 341778 268706 342334
rect 269262 341778 304706 342334
rect 305262 341778 340706 342334
rect 341262 341778 376706 342334
rect 377262 341778 412706 342334
rect 413262 341778 448706 342334
rect 449262 341778 484706 342334
rect 485262 341778 520706 342334
rect 521262 341778 556706 342334
rect 557262 341778 589182 342334
rect 589738 341778 592650 342334
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338058 -4854 338614
rect -4298 338058 12986 338614
rect 13542 338058 48986 338614
rect 49542 338058 84986 338614
rect 85542 338058 120986 338614
rect 121542 338058 156986 338614
rect 157542 338058 192986 338614
rect 193542 338058 228986 338614
rect 229542 338058 264986 338614
rect 265542 338058 300986 338614
rect 301542 338058 336986 338614
rect 337542 338058 372986 338614
rect 373542 338058 408986 338614
rect 409542 338058 444986 338614
rect 445542 338058 480986 338614
rect 481542 338058 516986 338614
rect 517542 338058 552986 338614
rect 553542 338058 588222 338614
rect 588778 338058 592650 338614
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334338 -3894 334894
rect -3338 334338 9266 334894
rect 9822 334338 45266 334894
rect 45822 334338 81266 334894
rect 81822 334338 117266 334894
rect 117822 334338 153266 334894
rect 153822 334338 189266 334894
rect 189822 334338 225266 334894
rect 225822 334338 261266 334894
rect 261822 334338 297266 334894
rect 297822 334338 333266 334894
rect 333822 334338 405266 334894
rect 405822 334338 441266 334894
rect 441822 334338 513266 334894
rect 513822 334338 549266 334894
rect 549822 334338 587262 334894
rect 587818 334338 592650 334894
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330618 -2934 331174
rect -2378 330618 5546 331174
rect 6102 330938 31610 331174
rect 31846 330938 41546 331174
rect 6102 330854 41546 330938
rect 6102 330618 31610 330854
rect 31846 330618 41546 330854
rect 42102 330938 62330 331174
rect 62566 330938 93050 331174
rect 93286 330938 113546 331174
rect 42102 330854 113546 330938
rect 42102 330618 62330 330854
rect 62566 330618 93050 330854
rect 93286 330618 113546 330854
rect 114102 330938 123770 331174
rect 124006 330938 149546 331174
rect 114102 330854 149546 330938
rect 114102 330618 123770 330854
rect 124006 330618 149546 330854
rect 150102 330938 154490 331174
rect 154726 330938 185210 331174
rect 185446 330938 215930 331174
rect 216166 330938 221546 331174
rect 150102 330854 221546 330938
rect 150102 330618 154490 330854
rect 154726 330618 185210 330854
rect 185446 330618 215930 330854
rect 216166 330618 221546 330854
rect 222102 330938 246650 331174
rect 246886 330938 257546 331174
rect 222102 330854 257546 330938
rect 222102 330618 246650 330854
rect 246886 330618 257546 330854
rect 258102 330938 277370 331174
rect 277606 330938 293546 331174
rect 258102 330854 293546 330938
rect 258102 330618 277370 330854
rect 277606 330618 293546 330854
rect 294102 330938 308090 331174
rect 308326 330938 329546 331174
rect 294102 330854 329546 330938
rect 294102 330618 308090 330854
rect 308326 330618 329546 330854
rect 330102 330938 338810 331174
rect 339046 330938 365546 331174
rect 330102 330854 365546 330938
rect 330102 330618 338810 330854
rect 339046 330618 365546 330854
rect 366102 330938 369530 331174
rect 369766 330938 400250 331174
rect 400486 330938 401546 331174
rect 366102 330854 401546 330938
rect 366102 330618 369530 330854
rect 369766 330618 400250 330854
rect 400486 330618 401546 330854
rect 402102 330938 430970 331174
rect 431206 330938 437546 331174
rect 402102 330854 437546 330938
rect 402102 330618 430970 330854
rect 431206 330618 437546 330854
rect 438102 330938 461690 331174
rect 461926 330938 473546 331174
rect 438102 330854 473546 330938
rect 438102 330618 461690 330854
rect 461926 330618 473546 330854
rect 474102 330938 492410 331174
rect 492646 330938 509546 331174
rect 474102 330854 509546 330938
rect 474102 330618 492410 330854
rect 492646 330618 509546 330854
rect 510102 330938 523130 331174
rect 523366 330938 545546 331174
rect 510102 330854 545546 330938
rect 510102 330618 523130 330854
rect 523366 330618 545546 330854
rect 546102 330938 553850 331174
rect 554086 330938 581546 331174
rect 546102 330854 581546 330938
rect 546102 330618 553850 330854
rect 554086 330618 581546 330854
rect 582102 330618 586302 331174
rect 586858 330618 592650 331174
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 326898 -1974 327454
rect -1418 326898 1826 327454
rect 2382 327218 16250 327454
rect 16486 327218 37826 327454
rect 2382 327134 37826 327218
rect 2382 326898 16250 327134
rect 16486 326898 37826 327134
rect 38382 327218 46970 327454
rect 47206 327218 73826 327454
rect 38382 327134 73826 327218
rect 38382 326898 46970 327134
rect 47206 326898 73826 327134
rect 74382 327218 77690 327454
rect 77926 327218 108410 327454
rect 108646 327218 109826 327454
rect 74382 327134 109826 327218
rect 74382 326898 77690 327134
rect 77926 326898 108410 327134
rect 108646 326898 109826 327134
rect 110382 327218 139130 327454
rect 139366 327218 145826 327454
rect 110382 327134 145826 327218
rect 110382 326898 139130 327134
rect 139366 326898 145826 327134
rect 146382 327218 169850 327454
rect 170086 327218 181826 327454
rect 146382 327134 181826 327218
rect 146382 326898 169850 327134
rect 170086 326898 181826 327134
rect 182382 327218 200570 327454
rect 200806 327218 217826 327454
rect 182382 327134 217826 327218
rect 182382 326898 200570 327134
rect 200806 326898 217826 327134
rect 218382 327218 231290 327454
rect 231526 327218 253826 327454
rect 218382 327134 253826 327218
rect 218382 326898 231290 327134
rect 231526 326898 253826 327134
rect 254382 327218 262010 327454
rect 262246 327218 289826 327454
rect 254382 327134 289826 327218
rect 254382 326898 262010 327134
rect 262246 326898 289826 327134
rect 290382 327218 292730 327454
rect 292966 327218 323450 327454
rect 323686 327218 325826 327454
rect 290382 327134 325826 327218
rect 290382 326898 292730 327134
rect 292966 326898 323450 327134
rect 323686 326898 325826 327134
rect 326382 327218 354170 327454
rect 354406 327218 361826 327454
rect 326382 327134 361826 327218
rect 326382 326898 354170 327134
rect 354406 326898 361826 327134
rect 362382 327218 384890 327454
rect 385126 327218 397826 327454
rect 362382 327134 397826 327218
rect 362382 326898 384890 327134
rect 385126 326898 397826 327134
rect 398382 327218 415610 327454
rect 415846 327218 433826 327454
rect 398382 327134 433826 327218
rect 398382 326898 415610 327134
rect 415846 326898 433826 327134
rect 434382 327218 446330 327454
rect 446566 327218 469826 327454
rect 434382 327134 469826 327218
rect 434382 326898 446330 327134
rect 446566 326898 469826 327134
rect 470382 327218 477050 327454
rect 477286 327218 505826 327454
rect 470382 327134 505826 327218
rect 470382 326898 477050 327134
rect 477286 326898 505826 327134
rect 506382 327218 507770 327454
rect 508006 327218 538490 327454
rect 538726 327218 541826 327454
rect 506382 327134 541826 327218
rect 506382 326898 507770 327134
rect 508006 326898 538490 327134
rect 538726 326898 541826 327134
rect 542382 327218 569210 327454
rect 569446 327218 577826 327454
rect 542382 327134 577826 327218
rect 542382 326898 569210 327134
rect 569446 326898 577826 327134
rect 578382 326898 585342 327454
rect 585898 326898 592650 327454
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 316938 -8694 317494
rect -8138 316938 27866 317494
rect 28422 316938 63866 317494
rect 64422 316938 99866 317494
rect 100422 316938 135866 317494
rect 136422 316938 171866 317494
rect 172422 316938 207866 317494
rect 208422 316938 243866 317494
rect 244422 316938 279866 317494
rect 280422 316938 315866 317494
rect 316422 316938 351866 317494
rect 352422 316938 387866 317494
rect 388422 316938 423866 317494
rect 424422 316938 459866 317494
rect 460422 316938 495866 317494
rect 496422 316938 531866 317494
rect 532422 316938 567866 317494
rect 568422 316938 592062 317494
rect 592618 316938 592650 317494
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313218 -7734 313774
rect -7178 313218 24146 313774
rect 24702 313218 60146 313774
rect 60702 313218 96146 313774
rect 96702 313218 132146 313774
rect 132702 313218 168146 313774
rect 168702 313218 204146 313774
rect 204702 313218 240146 313774
rect 240702 313218 276146 313774
rect 276702 313218 312146 313774
rect 312702 313218 348146 313774
rect 348702 313218 384146 313774
rect 384702 313218 420146 313774
rect 420702 313218 456146 313774
rect 456702 313218 528146 313774
rect 528702 313218 564146 313774
rect 564702 313218 591102 313774
rect 591658 313218 592650 313774
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309498 -6774 310054
rect -6218 309498 20426 310054
rect 20982 309498 56426 310054
rect 56982 309498 128426 310054
rect 128982 309498 164426 310054
rect 164982 309498 236426 310054
rect 236982 309498 272426 310054
rect 272982 309498 344426 310054
rect 344982 309498 380426 310054
rect 380982 309498 416426 310054
rect 416982 309498 452426 310054
rect 452982 309498 488426 310054
rect 488982 309498 524426 310054
rect 524982 309498 560426 310054
rect 560982 309498 590142 310054
rect 590698 309498 592650 310054
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 305778 -5814 306334
rect -5258 305778 16706 306334
rect 17262 305778 52706 306334
rect 53262 305778 88706 306334
rect 89262 305778 124706 306334
rect 125262 305778 160706 306334
rect 161262 305778 196706 306334
rect 197262 305778 232706 306334
rect 233262 305778 268706 306334
rect 269262 305778 304706 306334
rect 305262 305778 340706 306334
rect 341262 305778 376706 306334
rect 377262 305778 412706 306334
rect 413262 305778 448706 306334
rect 449262 305778 484706 306334
rect 485262 305778 520706 306334
rect 521262 305778 556706 306334
rect 557262 305778 589182 306334
rect 589738 305778 592650 306334
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302058 -4854 302614
rect -4298 302058 12986 302614
rect 13542 302058 48986 302614
rect 49542 302058 84986 302614
rect 85542 302058 120986 302614
rect 121542 302058 156986 302614
rect 157542 302058 192986 302614
rect 193542 302058 228986 302614
rect 229542 302058 264986 302614
rect 265542 302058 300986 302614
rect 301542 302058 336986 302614
rect 337542 302058 372986 302614
rect 373542 302058 408986 302614
rect 409542 302058 444986 302614
rect 445542 302058 480986 302614
rect 481542 302058 516986 302614
rect 517542 302058 552986 302614
rect 553542 302058 588222 302614
rect 588778 302058 592650 302614
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298338 -3894 298894
rect -3338 298338 9266 298894
rect 9822 298338 45266 298894
rect 45822 298338 81266 298894
rect 81822 298338 117266 298894
rect 117822 298338 153266 298894
rect 153822 298338 189266 298894
rect 189822 298338 225266 298894
rect 225822 298338 261266 298894
rect 261822 298338 297266 298894
rect 297822 298338 333266 298894
rect 333822 298338 405266 298894
rect 405822 298338 441266 298894
rect 441822 298338 513266 298894
rect 513822 298338 549266 298894
rect 549822 298338 587262 298894
rect 587818 298338 592650 298894
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294618 -2934 295174
rect -2378 294618 5546 295174
rect 6102 294938 31610 295174
rect 31846 294938 41546 295174
rect 6102 294854 41546 294938
rect 6102 294618 31610 294854
rect 31846 294618 41546 294854
rect 42102 294938 62330 295174
rect 62566 294938 93050 295174
rect 93286 294938 113546 295174
rect 42102 294854 113546 294938
rect 42102 294618 62330 294854
rect 62566 294618 93050 294854
rect 93286 294618 113546 294854
rect 114102 294938 123770 295174
rect 124006 294938 149546 295174
rect 114102 294854 149546 294938
rect 114102 294618 123770 294854
rect 124006 294618 149546 294854
rect 150102 294938 154490 295174
rect 154726 294938 185210 295174
rect 185446 294938 215930 295174
rect 216166 294938 221546 295174
rect 150102 294854 221546 294938
rect 150102 294618 154490 294854
rect 154726 294618 185210 294854
rect 185446 294618 215930 294854
rect 216166 294618 221546 294854
rect 222102 294938 246650 295174
rect 246886 294938 257546 295174
rect 222102 294854 257546 294938
rect 222102 294618 246650 294854
rect 246886 294618 257546 294854
rect 258102 294938 277370 295174
rect 277606 294938 293546 295174
rect 258102 294854 293546 294938
rect 258102 294618 277370 294854
rect 277606 294618 293546 294854
rect 294102 294938 308090 295174
rect 308326 294938 329546 295174
rect 294102 294854 329546 294938
rect 294102 294618 308090 294854
rect 308326 294618 329546 294854
rect 330102 294938 338810 295174
rect 339046 294938 365546 295174
rect 330102 294854 365546 294938
rect 330102 294618 338810 294854
rect 339046 294618 365546 294854
rect 366102 294938 369530 295174
rect 369766 294938 400250 295174
rect 400486 294938 401546 295174
rect 366102 294854 401546 294938
rect 366102 294618 369530 294854
rect 369766 294618 400250 294854
rect 400486 294618 401546 294854
rect 402102 294938 430970 295174
rect 431206 294938 437546 295174
rect 402102 294854 437546 294938
rect 402102 294618 430970 294854
rect 431206 294618 437546 294854
rect 438102 294938 461690 295174
rect 461926 294938 473546 295174
rect 438102 294854 473546 294938
rect 438102 294618 461690 294854
rect 461926 294618 473546 294854
rect 474102 294938 492410 295174
rect 492646 294938 509546 295174
rect 474102 294854 509546 294938
rect 474102 294618 492410 294854
rect 492646 294618 509546 294854
rect 510102 294938 523130 295174
rect 523366 294938 545546 295174
rect 510102 294854 545546 294938
rect 510102 294618 523130 294854
rect 523366 294618 545546 294854
rect 546102 294938 553850 295174
rect 554086 294938 581546 295174
rect 546102 294854 581546 294938
rect 546102 294618 553850 294854
rect 554086 294618 581546 294854
rect 582102 294618 586302 295174
rect 586858 294618 592650 295174
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 290898 -1974 291454
rect -1418 290898 1826 291454
rect 2382 291218 16250 291454
rect 16486 291218 37826 291454
rect 2382 291134 37826 291218
rect 2382 290898 16250 291134
rect 16486 290898 37826 291134
rect 38382 291218 46970 291454
rect 47206 291218 73826 291454
rect 38382 291134 73826 291218
rect 38382 290898 46970 291134
rect 47206 290898 73826 291134
rect 74382 291218 77690 291454
rect 77926 291218 108410 291454
rect 108646 291218 109826 291454
rect 74382 291134 109826 291218
rect 74382 290898 77690 291134
rect 77926 290898 108410 291134
rect 108646 290898 109826 291134
rect 110382 291218 139130 291454
rect 139366 291218 145826 291454
rect 110382 291134 145826 291218
rect 110382 290898 139130 291134
rect 139366 290898 145826 291134
rect 146382 291218 169850 291454
rect 170086 291218 181826 291454
rect 146382 291134 181826 291218
rect 146382 290898 169850 291134
rect 170086 290898 181826 291134
rect 182382 291218 200570 291454
rect 200806 291218 217826 291454
rect 182382 291134 217826 291218
rect 182382 290898 200570 291134
rect 200806 290898 217826 291134
rect 218382 291218 231290 291454
rect 231526 291218 253826 291454
rect 218382 291134 253826 291218
rect 218382 290898 231290 291134
rect 231526 290898 253826 291134
rect 254382 291218 262010 291454
rect 262246 291218 289826 291454
rect 254382 291134 289826 291218
rect 254382 290898 262010 291134
rect 262246 290898 289826 291134
rect 290382 291218 292730 291454
rect 292966 291218 323450 291454
rect 323686 291218 325826 291454
rect 290382 291134 325826 291218
rect 290382 290898 292730 291134
rect 292966 290898 323450 291134
rect 323686 290898 325826 291134
rect 326382 291218 354170 291454
rect 354406 291218 361826 291454
rect 326382 291134 361826 291218
rect 326382 290898 354170 291134
rect 354406 290898 361826 291134
rect 362382 291218 384890 291454
rect 385126 291218 397826 291454
rect 362382 291134 397826 291218
rect 362382 290898 384890 291134
rect 385126 290898 397826 291134
rect 398382 291218 415610 291454
rect 415846 291218 433826 291454
rect 398382 291134 433826 291218
rect 398382 290898 415610 291134
rect 415846 290898 433826 291134
rect 434382 291218 446330 291454
rect 446566 291218 469826 291454
rect 434382 291134 469826 291218
rect 434382 290898 446330 291134
rect 446566 290898 469826 291134
rect 470382 291218 477050 291454
rect 477286 291218 505826 291454
rect 470382 291134 505826 291218
rect 470382 290898 477050 291134
rect 477286 290898 505826 291134
rect 506382 291218 507770 291454
rect 508006 291218 538490 291454
rect 538726 291218 541826 291454
rect 506382 291134 541826 291218
rect 506382 290898 507770 291134
rect 508006 290898 538490 291134
rect 538726 290898 541826 291134
rect 542382 291218 569210 291454
rect 569446 291218 577826 291454
rect 542382 291134 577826 291218
rect 542382 290898 569210 291134
rect 569446 290898 577826 291134
rect 578382 290898 585342 291454
rect 585898 290898 592650 291454
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 280938 -8694 281494
rect -8138 280938 27866 281494
rect 28422 280938 63866 281494
rect 64422 280938 99866 281494
rect 100422 280938 135866 281494
rect 136422 280938 171866 281494
rect 172422 280938 207866 281494
rect 208422 280938 243866 281494
rect 244422 280938 279866 281494
rect 280422 280938 315866 281494
rect 316422 280938 351866 281494
rect 352422 280938 387866 281494
rect 388422 280938 423866 281494
rect 424422 280938 459866 281494
rect 460422 280938 495866 281494
rect 496422 280938 531866 281494
rect 532422 280938 567866 281494
rect 568422 280938 592062 281494
rect 592618 280938 592650 281494
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277218 -7734 277774
rect -7178 277218 24146 277774
rect 24702 277218 60146 277774
rect 60702 277218 96146 277774
rect 96702 277218 132146 277774
rect 132702 277218 168146 277774
rect 168702 277218 204146 277774
rect 204702 277218 240146 277774
rect 240702 277218 276146 277774
rect 276702 277218 312146 277774
rect 312702 277218 348146 277774
rect 348702 277218 384146 277774
rect 384702 277218 420146 277774
rect 420702 277218 456146 277774
rect 456702 277218 528146 277774
rect 528702 277218 564146 277774
rect 564702 277218 591102 277774
rect 591658 277218 592650 277774
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273498 -6774 274054
rect -6218 273498 20426 274054
rect 20982 273498 56426 274054
rect 56982 273498 128426 274054
rect 128982 273498 164426 274054
rect 164982 273498 236426 274054
rect 236982 273498 272426 274054
rect 272982 273498 344426 274054
rect 344982 273498 380426 274054
rect 380982 273498 416426 274054
rect 416982 273498 452426 274054
rect 452982 273498 488426 274054
rect 488982 273498 524426 274054
rect 524982 273498 560426 274054
rect 560982 273498 590142 274054
rect 590698 273498 592650 274054
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 269778 -5814 270334
rect -5258 269778 16706 270334
rect 17262 269778 52706 270334
rect 53262 269778 88706 270334
rect 89262 269778 124706 270334
rect 125262 269778 160706 270334
rect 161262 269778 196706 270334
rect 197262 269778 232706 270334
rect 233262 269778 268706 270334
rect 269262 269778 304706 270334
rect 305262 269778 340706 270334
rect 341262 269778 376706 270334
rect 377262 269778 412706 270334
rect 413262 269778 448706 270334
rect 449262 269778 484706 270334
rect 485262 269778 520706 270334
rect 521262 269778 556706 270334
rect 557262 269778 589182 270334
rect 589738 269778 592650 270334
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266058 -4854 266614
rect -4298 266058 12986 266614
rect 13542 266058 48986 266614
rect 49542 266058 84986 266614
rect 85542 266058 120986 266614
rect 121542 266058 156986 266614
rect 157542 266058 192986 266614
rect 193542 266058 228986 266614
rect 229542 266058 264986 266614
rect 265542 266058 300986 266614
rect 301542 266058 336986 266614
rect 337542 266058 372986 266614
rect 373542 266058 408986 266614
rect 409542 266058 444986 266614
rect 445542 266058 480986 266614
rect 481542 266058 516986 266614
rect 517542 266058 552986 266614
rect 553542 266058 588222 266614
rect 588778 266058 592650 266614
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262338 -3894 262894
rect -3338 262338 9266 262894
rect 9822 262338 45266 262894
rect 45822 262338 81266 262894
rect 81822 262338 117266 262894
rect 117822 262338 153266 262894
rect 153822 262338 189266 262894
rect 189822 262338 225266 262894
rect 225822 262338 261266 262894
rect 261822 262338 297266 262894
rect 297822 262338 333266 262894
rect 333822 262338 405266 262894
rect 405822 262338 441266 262894
rect 441822 262338 513266 262894
rect 513822 262338 549266 262894
rect 549822 262338 587262 262894
rect 587818 262338 592650 262894
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258618 -2934 259174
rect -2378 258618 5546 259174
rect 6102 258938 31610 259174
rect 31846 258938 41546 259174
rect 6102 258854 41546 258938
rect 6102 258618 31610 258854
rect 31846 258618 41546 258854
rect 42102 258938 62330 259174
rect 62566 258938 93050 259174
rect 93286 258938 113546 259174
rect 42102 258854 113546 258938
rect 42102 258618 62330 258854
rect 62566 258618 93050 258854
rect 93286 258618 113546 258854
rect 114102 258938 123770 259174
rect 124006 258938 149546 259174
rect 114102 258854 149546 258938
rect 114102 258618 123770 258854
rect 124006 258618 149546 258854
rect 150102 258938 154490 259174
rect 154726 258938 185210 259174
rect 185446 258938 215930 259174
rect 216166 258938 221546 259174
rect 150102 258854 221546 258938
rect 150102 258618 154490 258854
rect 154726 258618 185210 258854
rect 185446 258618 215930 258854
rect 216166 258618 221546 258854
rect 222102 258938 246650 259174
rect 246886 258938 257546 259174
rect 222102 258854 257546 258938
rect 222102 258618 246650 258854
rect 246886 258618 257546 258854
rect 258102 258938 277370 259174
rect 277606 258938 293546 259174
rect 258102 258854 293546 258938
rect 258102 258618 277370 258854
rect 277606 258618 293546 258854
rect 294102 258938 308090 259174
rect 308326 258938 329546 259174
rect 294102 258854 329546 258938
rect 294102 258618 308090 258854
rect 308326 258618 329546 258854
rect 330102 258938 338810 259174
rect 339046 258938 365546 259174
rect 330102 258854 365546 258938
rect 330102 258618 338810 258854
rect 339046 258618 365546 258854
rect 366102 258938 369530 259174
rect 369766 258938 400250 259174
rect 400486 258938 401546 259174
rect 366102 258854 401546 258938
rect 366102 258618 369530 258854
rect 369766 258618 400250 258854
rect 400486 258618 401546 258854
rect 402102 258938 430970 259174
rect 431206 258938 437546 259174
rect 402102 258854 437546 258938
rect 402102 258618 430970 258854
rect 431206 258618 437546 258854
rect 438102 258938 461690 259174
rect 461926 258938 473546 259174
rect 438102 258854 473546 258938
rect 438102 258618 461690 258854
rect 461926 258618 473546 258854
rect 474102 258938 492410 259174
rect 492646 258938 509546 259174
rect 474102 258854 509546 258938
rect 474102 258618 492410 258854
rect 492646 258618 509546 258854
rect 510102 258938 523130 259174
rect 523366 258938 545546 259174
rect 510102 258854 545546 258938
rect 510102 258618 523130 258854
rect 523366 258618 545546 258854
rect 546102 258938 553850 259174
rect 554086 258938 581546 259174
rect 546102 258854 581546 258938
rect 546102 258618 553850 258854
rect 554086 258618 581546 258854
rect 582102 258618 586302 259174
rect 586858 258618 592650 259174
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 254898 -1974 255454
rect -1418 254898 1826 255454
rect 2382 255218 16250 255454
rect 16486 255218 37826 255454
rect 2382 255134 37826 255218
rect 2382 254898 16250 255134
rect 16486 254898 37826 255134
rect 38382 255218 46970 255454
rect 47206 255218 73826 255454
rect 38382 255134 73826 255218
rect 38382 254898 46970 255134
rect 47206 254898 73826 255134
rect 74382 255218 77690 255454
rect 77926 255218 108410 255454
rect 108646 255218 109826 255454
rect 74382 255134 109826 255218
rect 74382 254898 77690 255134
rect 77926 254898 108410 255134
rect 108646 254898 109826 255134
rect 110382 255218 139130 255454
rect 139366 255218 145826 255454
rect 110382 255134 145826 255218
rect 110382 254898 139130 255134
rect 139366 254898 145826 255134
rect 146382 255218 169850 255454
rect 170086 255218 181826 255454
rect 146382 255134 181826 255218
rect 146382 254898 169850 255134
rect 170086 254898 181826 255134
rect 182382 255218 200570 255454
rect 200806 255218 217826 255454
rect 182382 255134 217826 255218
rect 182382 254898 200570 255134
rect 200806 254898 217826 255134
rect 218382 255218 231290 255454
rect 231526 255218 253826 255454
rect 218382 255134 253826 255218
rect 218382 254898 231290 255134
rect 231526 254898 253826 255134
rect 254382 255218 262010 255454
rect 262246 255218 289826 255454
rect 254382 255134 289826 255218
rect 254382 254898 262010 255134
rect 262246 254898 289826 255134
rect 290382 255218 292730 255454
rect 292966 255218 323450 255454
rect 323686 255218 325826 255454
rect 290382 255134 325826 255218
rect 290382 254898 292730 255134
rect 292966 254898 323450 255134
rect 323686 254898 325826 255134
rect 326382 255218 354170 255454
rect 354406 255218 361826 255454
rect 326382 255134 361826 255218
rect 326382 254898 354170 255134
rect 354406 254898 361826 255134
rect 362382 255218 384890 255454
rect 385126 255218 397826 255454
rect 362382 255134 397826 255218
rect 362382 254898 384890 255134
rect 385126 254898 397826 255134
rect 398382 255218 415610 255454
rect 415846 255218 433826 255454
rect 398382 255134 433826 255218
rect 398382 254898 415610 255134
rect 415846 254898 433826 255134
rect 434382 255218 446330 255454
rect 446566 255218 469826 255454
rect 434382 255134 469826 255218
rect 434382 254898 446330 255134
rect 446566 254898 469826 255134
rect 470382 255218 477050 255454
rect 477286 255218 505826 255454
rect 470382 255134 505826 255218
rect 470382 254898 477050 255134
rect 477286 254898 505826 255134
rect 506382 255218 507770 255454
rect 508006 255218 538490 255454
rect 538726 255218 541826 255454
rect 506382 255134 541826 255218
rect 506382 254898 507770 255134
rect 508006 254898 538490 255134
rect 538726 254898 541826 255134
rect 542382 255218 569210 255454
rect 569446 255218 577826 255454
rect 542382 255134 577826 255218
rect 542382 254898 569210 255134
rect 569446 254898 577826 255134
rect 578382 254898 585342 255454
rect 585898 254898 592650 255454
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 244938 -8694 245494
rect -8138 244938 27866 245494
rect 28422 244938 63866 245494
rect 64422 244938 99866 245494
rect 100422 244938 135866 245494
rect 136422 244938 171866 245494
rect 172422 244938 207866 245494
rect 208422 244938 243866 245494
rect 244422 244938 279866 245494
rect 280422 244938 315866 245494
rect 316422 244938 351866 245494
rect 352422 244938 387866 245494
rect 388422 244938 423866 245494
rect 424422 244938 459866 245494
rect 460422 244938 495866 245494
rect 496422 244938 531866 245494
rect 532422 244938 567866 245494
rect 568422 244938 592062 245494
rect 592618 244938 592650 245494
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241218 -7734 241774
rect -7178 241218 24146 241774
rect 24702 241218 60146 241774
rect 60702 241218 96146 241774
rect 96702 241218 132146 241774
rect 132702 241218 168146 241774
rect 168702 241218 204146 241774
rect 204702 241218 240146 241774
rect 240702 241218 276146 241774
rect 276702 241218 312146 241774
rect 312702 241218 348146 241774
rect 348702 241218 384146 241774
rect 384702 241218 420146 241774
rect 420702 241218 456146 241774
rect 456702 241218 528146 241774
rect 528702 241218 564146 241774
rect 564702 241218 591102 241774
rect 591658 241218 592650 241774
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237498 -6774 238054
rect -6218 237498 20426 238054
rect 20982 237498 56426 238054
rect 56982 237498 128426 238054
rect 128982 237498 164426 238054
rect 164982 237498 236426 238054
rect 236982 237498 272426 238054
rect 272982 237498 344426 238054
rect 344982 237498 380426 238054
rect 380982 237498 416426 238054
rect 416982 237498 452426 238054
rect 452982 237498 488426 238054
rect 488982 237498 524426 238054
rect 524982 237498 560426 238054
rect 560982 237498 590142 238054
rect 590698 237498 592650 238054
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 233778 -5814 234334
rect -5258 233778 16706 234334
rect 17262 233778 52706 234334
rect 53262 233778 88706 234334
rect 89262 233778 124706 234334
rect 125262 233778 160706 234334
rect 161262 233778 196706 234334
rect 197262 233778 232706 234334
rect 233262 233778 268706 234334
rect 269262 233778 304706 234334
rect 305262 233778 340706 234334
rect 341262 233778 376706 234334
rect 377262 233778 412706 234334
rect 413262 233778 448706 234334
rect 449262 233778 484706 234334
rect 485262 233778 520706 234334
rect 521262 233778 556706 234334
rect 557262 233778 589182 234334
rect 589738 233778 592650 234334
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230058 -4854 230614
rect -4298 230058 12986 230614
rect 13542 230058 48986 230614
rect 49542 230058 84986 230614
rect 85542 230058 120986 230614
rect 121542 230058 156986 230614
rect 157542 230058 192986 230614
rect 193542 230058 228986 230614
rect 229542 230058 264986 230614
rect 265542 230058 300986 230614
rect 301542 230058 336986 230614
rect 337542 230058 372986 230614
rect 373542 230058 408986 230614
rect 409542 230058 444986 230614
rect 445542 230058 480986 230614
rect 481542 230058 516986 230614
rect 517542 230058 552986 230614
rect 553542 230058 588222 230614
rect 588778 230058 592650 230614
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226338 -3894 226894
rect -3338 226338 9266 226894
rect 9822 226338 45266 226894
rect 45822 226338 81266 226894
rect 81822 226338 117266 226894
rect 117822 226338 153266 226894
rect 153822 226338 189266 226894
rect 189822 226338 225266 226894
rect 225822 226338 261266 226894
rect 261822 226338 297266 226894
rect 297822 226338 333266 226894
rect 333822 226338 405266 226894
rect 405822 226338 441266 226894
rect 441822 226338 513266 226894
rect 513822 226338 549266 226894
rect 549822 226338 587262 226894
rect 587818 226338 592650 226894
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222618 -2934 223174
rect -2378 222618 5546 223174
rect 6102 222938 31610 223174
rect 31846 222938 41546 223174
rect 6102 222854 41546 222938
rect 6102 222618 31610 222854
rect 31846 222618 41546 222854
rect 42102 222938 62330 223174
rect 62566 222938 93050 223174
rect 93286 222938 113546 223174
rect 42102 222854 113546 222938
rect 42102 222618 62330 222854
rect 62566 222618 93050 222854
rect 93286 222618 113546 222854
rect 114102 222938 123770 223174
rect 124006 222938 149546 223174
rect 114102 222854 149546 222938
rect 114102 222618 123770 222854
rect 124006 222618 149546 222854
rect 150102 222938 154490 223174
rect 154726 222938 185210 223174
rect 185446 222938 215930 223174
rect 216166 222938 221546 223174
rect 150102 222854 221546 222938
rect 150102 222618 154490 222854
rect 154726 222618 185210 222854
rect 185446 222618 215930 222854
rect 216166 222618 221546 222854
rect 222102 222938 246650 223174
rect 246886 222938 257546 223174
rect 222102 222854 257546 222938
rect 222102 222618 246650 222854
rect 246886 222618 257546 222854
rect 258102 222938 277370 223174
rect 277606 222938 293546 223174
rect 258102 222854 293546 222938
rect 258102 222618 277370 222854
rect 277606 222618 293546 222854
rect 294102 222938 308090 223174
rect 308326 222938 329546 223174
rect 294102 222854 329546 222938
rect 294102 222618 308090 222854
rect 308326 222618 329546 222854
rect 330102 222938 338810 223174
rect 339046 222938 365546 223174
rect 330102 222854 365546 222938
rect 330102 222618 338810 222854
rect 339046 222618 365546 222854
rect 366102 222938 369530 223174
rect 369766 222938 400250 223174
rect 400486 222938 401546 223174
rect 366102 222854 401546 222938
rect 366102 222618 369530 222854
rect 369766 222618 400250 222854
rect 400486 222618 401546 222854
rect 402102 222938 430970 223174
rect 431206 222938 437546 223174
rect 402102 222854 437546 222938
rect 402102 222618 430970 222854
rect 431206 222618 437546 222854
rect 438102 222938 461690 223174
rect 461926 222938 473546 223174
rect 438102 222854 473546 222938
rect 438102 222618 461690 222854
rect 461926 222618 473546 222854
rect 474102 222938 492410 223174
rect 492646 222938 509546 223174
rect 474102 222854 509546 222938
rect 474102 222618 492410 222854
rect 492646 222618 509546 222854
rect 510102 222938 523130 223174
rect 523366 222938 545546 223174
rect 510102 222854 545546 222938
rect 510102 222618 523130 222854
rect 523366 222618 545546 222854
rect 546102 222938 553850 223174
rect 554086 222938 581546 223174
rect 546102 222854 581546 222938
rect 546102 222618 553850 222854
rect 554086 222618 581546 222854
rect 582102 222618 586302 223174
rect 586858 222618 592650 223174
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 218898 -1974 219454
rect -1418 218898 1826 219454
rect 2382 219218 16250 219454
rect 16486 219218 37826 219454
rect 2382 219134 37826 219218
rect 2382 218898 16250 219134
rect 16486 218898 37826 219134
rect 38382 219218 46970 219454
rect 47206 219218 73826 219454
rect 38382 219134 73826 219218
rect 38382 218898 46970 219134
rect 47206 218898 73826 219134
rect 74382 219218 77690 219454
rect 77926 219218 108410 219454
rect 108646 219218 109826 219454
rect 74382 219134 109826 219218
rect 74382 218898 77690 219134
rect 77926 218898 108410 219134
rect 108646 218898 109826 219134
rect 110382 219218 139130 219454
rect 139366 219218 145826 219454
rect 110382 219134 145826 219218
rect 110382 218898 139130 219134
rect 139366 218898 145826 219134
rect 146382 219218 169850 219454
rect 170086 219218 181826 219454
rect 146382 219134 181826 219218
rect 146382 218898 169850 219134
rect 170086 218898 181826 219134
rect 182382 219218 200570 219454
rect 200806 219218 217826 219454
rect 182382 219134 217826 219218
rect 182382 218898 200570 219134
rect 200806 218898 217826 219134
rect 218382 219218 231290 219454
rect 231526 219218 253826 219454
rect 218382 219134 253826 219218
rect 218382 218898 231290 219134
rect 231526 218898 253826 219134
rect 254382 219218 262010 219454
rect 262246 219218 289826 219454
rect 254382 219134 289826 219218
rect 254382 218898 262010 219134
rect 262246 218898 289826 219134
rect 290382 219218 292730 219454
rect 292966 219218 323450 219454
rect 323686 219218 325826 219454
rect 290382 219134 325826 219218
rect 290382 218898 292730 219134
rect 292966 218898 323450 219134
rect 323686 218898 325826 219134
rect 326382 219218 354170 219454
rect 354406 219218 361826 219454
rect 326382 219134 361826 219218
rect 326382 218898 354170 219134
rect 354406 218898 361826 219134
rect 362382 219218 384890 219454
rect 385126 219218 397826 219454
rect 362382 219134 397826 219218
rect 362382 218898 384890 219134
rect 385126 218898 397826 219134
rect 398382 219218 415610 219454
rect 415846 219218 433826 219454
rect 398382 219134 433826 219218
rect 398382 218898 415610 219134
rect 415846 218898 433826 219134
rect 434382 219218 446330 219454
rect 446566 219218 469826 219454
rect 434382 219134 469826 219218
rect 434382 218898 446330 219134
rect 446566 218898 469826 219134
rect 470382 219218 477050 219454
rect 477286 219218 505826 219454
rect 470382 219134 505826 219218
rect 470382 218898 477050 219134
rect 477286 218898 505826 219134
rect 506382 219218 507770 219454
rect 508006 219218 538490 219454
rect 538726 219218 541826 219454
rect 506382 219134 541826 219218
rect 506382 218898 507770 219134
rect 508006 218898 538490 219134
rect 538726 218898 541826 219134
rect 542382 219218 569210 219454
rect 569446 219218 577826 219454
rect 542382 219134 577826 219218
rect 542382 218898 569210 219134
rect 569446 218898 577826 219134
rect 578382 218898 585342 219454
rect 585898 218898 592650 219454
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 208938 -8694 209494
rect -8138 208938 27866 209494
rect 28422 208938 63866 209494
rect 64422 208938 99866 209494
rect 100422 208938 135866 209494
rect 136422 208938 171866 209494
rect 172422 208938 207866 209494
rect 208422 208938 243866 209494
rect 244422 208938 279866 209494
rect 280422 208938 315866 209494
rect 316422 208938 351866 209494
rect 352422 208938 387866 209494
rect 388422 208938 423866 209494
rect 424422 208938 459866 209494
rect 460422 208938 495866 209494
rect 496422 208938 531866 209494
rect 532422 208938 567866 209494
rect 568422 208938 592062 209494
rect 592618 208938 592650 209494
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205218 -7734 205774
rect -7178 205218 24146 205774
rect 24702 205218 60146 205774
rect 60702 205218 96146 205774
rect 96702 205218 132146 205774
rect 132702 205218 168146 205774
rect 168702 205218 204146 205774
rect 204702 205218 240146 205774
rect 240702 205218 276146 205774
rect 276702 205218 312146 205774
rect 312702 205218 348146 205774
rect 348702 205218 384146 205774
rect 384702 205218 420146 205774
rect 420702 205218 456146 205774
rect 456702 205218 528146 205774
rect 528702 205218 564146 205774
rect 564702 205218 591102 205774
rect 591658 205218 592650 205774
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201498 -6774 202054
rect -6218 201498 20426 202054
rect 20982 201498 56426 202054
rect 56982 201498 128426 202054
rect 128982 201498 164426 202054
rect 164982 201498 236426 202054
rect 236982 201498 272426 202054
rect 272982 201498 344426 202054
rect 344982 201498 380426 202054
rect 380982 201498 416426 202054
rect 416982 201498 452426 202054
rect 452982 201498 488426 202054
rect 488982 201498 524426 202054
rect 524982 201498 560426 202054
rect 560982 201498 590142 202054
rect 590698 201498 592650 202054
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 197778 -5814 198334
rect -5258 197778 16706 198334
rect 17262 197778 52706 198334
rect 53262 197778 88706 198334
rect 89262 197778 124706 198334
rect 125262 197778 160706 198334
rect 161262 197778 196706 198334
rect 197262 197778 232706 198334
rect 233262 197778 268706 198334
rect 269262 197778 304706 198334
rect 305262 197778 340706 198334
rect 341262 197778 376706 198334
rect 377262 197778 412706 198334
rect 413262 197778 448706 198334
rect 449262 197778 484706 198334
rect 485262 197778 520706 198334
rect 521262 197778 556706 198334
rect 557262 197778 589182 198334
rect 589738 197778 592650 198334
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194058 -4854 194614
rect -4298 194058 12986 194614
rect 13542 194058 48986 194614
rect 49542 194058 84986 194614
rect 85542 194058 120986 194614
rect 121542 194058 156986 194614
rect 157542 194058 192986 194614
rect 193542 194058 228986 194614
rect 229542 194058 264986 194614
rect 265542 194058 300986 194614
rect 301542 194058 336986 194614
rect 337542 194058 372986 194614
rect 373542 194058 408986 194614
rect 409542 194058 444986 194614
rect 445542 194058 480986 194614
rect 481542 194058 516986 194614
rect 517542 194058 552986 194614
rect 553542 194058 588222 194614
rect 588778 194058 592650 194614
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190338 -3894 190894
rect -3338 190338 9266 190894
rect 9822 190338 45266 190894
rect 45822 190338 81266 190894
rect 81822 190338 117266 190894
rect 117822 190338 153266 190894
rect 153822 190338 189266 190894
rect 189822 190338 225266 190894
rect 225822 190338 261266 190894
rect 261822 190338 297266 190894
rect 297822 190338 333266 190894
rect 333822 190338 405266 190894
rect 405822 190338 441266 190894
rect 441822 190338 513266 190894
rect 513822 190338 549266 190894
rect 549822 190338 587262 190894
rect 587818 190338 592650 190894
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186618 -2934 187174
rect -2378 186618 5546 187174
rect 6102 186938 31610 187174
rect 31846 186938 41546 187174
rect 6102 186854 41546 186938
rect 6102 186618 31610 186854
rect 31846 186618 41546 186854
rect 42102 186938 62330 187174
rect 62566 186938 93050 187174
rect 93286 186938 113546 187174
rect 42102 186854 113546 186938
rect 42102 186618 62330 186854
rect 62566 186618 93050 186854
rect 93286 186618 113546 186854
rect 114102 186938 123770 187174
rect 124006 186938 149546 187174
rect 114102 186854 149546 186938
rect 114102 186618 123770 186854
rect 124006 186618 149546 186854
rect 150102 186938 154490 187174
rect 154726 186938 185210 187174
rect 185446 186938 215930 187174
rect 216166 186938 221546 187174
rect 150102 186854 221546 186938
rect 150102 186618 154490 186854
rect 154726 186618 185210 186854
rect 185446 186618 215930 186854
rect 216166 186618 221546 186854
rect 222102 186938 246650 187174
rect 246886 186938 257546 187174
rect 222102 186854 257546 186938
rect 222102 186618 246650 186854
rect 246886 186618 257546 186854
rect 258102 186938 277370 187174
rect 277606 186938 293546 187174
rect 258102 186854 293546 186938
rect 258102 186618 277370 186854
rect 277606 186618 293546 186854
rect 294102 186938 308090 187174
rect 308326 186938 329546 187174
rect 294102 186854 329546 186938
rect 294102 186618 308090 186854
rect 308326 186618 329546 186854
rect 330102 186938 338810 187174
rect 339046 186938 365546 187174
rect 330102 186854 365546 186938
rect 330102 186618 338810 186854
rect 339046 186618 365546 186854
rect 366102 186938 369530 187174
rect 369766 186938 400250 187174
rect 400486 186938 401546 187174
rect 366102 186854 401546 186938
rect 366102 186618 369530 186854
rect 369766 186618 400250 186854
rect 400486 186618 401546 186854
rect 402102 186938 430970 187174
rect 431206 186938 437546 187174
rect 402102 186854 437546 186938
rect 402102 186618 430970 186854
rect 431206 186618 437546 186854
rect 438102 186938 461690 187174
rect 461926 186938 473546 187174
rect 438102 186854 473546 186938
rect 438102 186618 461690 186854
rect 461926 186618 473546 186854
rect 474102 186938 492410 187174
rect 492646 186938 509546 187174
rect 474102 186854 509546 186938
rect 474102 186618 492410 186854
rect 492646 186618 509546 186854
rect 510102 186938 523130 187174
rect 523366 186938 545546 187174
rect 510102 186854 545546 186938
rect 510102 186618 523130 186854
rect 523366 186618 545546 186854
rect 546102 186938 553850 187174
rect 554086 186938 581546 187174
rect 546102 186854 581546 186938
rect 546102 186618 553850 186854
rect 554086 186618 581546 186854
rect 582102 186618 586302 187174
rect 586858 186618 592650 187174
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 182898 -1974 183454
rect -1418 182898 1826 183454
rect 2382 183218 16250 183454
rect 16486 183218 37826 183454
rect 2382 183134 37826 183218
rect 2382 182898 16250 183134
rect 16486 182898 37826 183134
rect 38382 183218 46970 183454
rect 47206 183218 73826 183454
rect 38382 183134 73826 183218
rect 38382 182898 46970 183134
rect 47206 182898 73826 183134
rect 74382 183218 77690 183454
rect 77926 183218 108410 183454
rect 108646 183218 109826 183454
rect 74382 183134 109826 183218
rect 74382 182898 77690 183134
rect 77926 182898 108410 183134
rect 108646 182898 109826 183134
rect 110382 183218 139130 183454
rect 139366 183218 145826 183454
rect 110382 183134 145826 183218
rect 110382 182898 139130 183134
rect 139366 182898 145826 183134
rect 146382 183218 169850 183454
rect 170086 183218 181826 183454
rect 146382 183134 181826 183218
rect 146382 182898 169850 183134
rect 170086 182898 181826 183134
rect 182382 183218 200570 183454
rect 200806 183218 217826 183454
rect 182382 183134 217826 183218
rect 182382 182898 200570 183134
rect 200806 182898 217826 183134
rect 218382 183218 231290 183454
rect 231526 183218 253826 183454
rect 218382 183134 253826 183218
rect 218382 182898 231290 183134
rect 231526 182898 253826 183134
rect 254382 183218 262010 183454
rect 262246 183218 289826 183454
rect 254382 183134 289826 183218
rect 254382 182898 262010 183134
rect 262246 182898 289826 183134
rect 290382 183218 292730 183454
rect 292966 183218 323450 183454
rect 323686 183218 325826 183454
rect 290382 183134 325826 183218
rect 290382 182898 292730 183134
rect 292966 182898 323450 183134
rect 323686 182898 325826 183134
rect 326382 183218 354170 183454
rect 354406 183218 361826 183454
rect 326382 183134 361826 183218
rect 326382 182898 354170 183134
rect 354406 182898 361826 183134
rect 362382 183218 384890 183454
rect 385126 183218 397826 183454
rect 362382 183134 397826 183218
rect 362382 182898 384890 183134
rect 385126 182898 397826 183134
rect 398382 183218 415610 183454
rect 415846 183218 433826 183454
rect 398382 183134 433826 183218
rect 398382 182898 415610 183134
rect 415846 182898 433826 183134
rect 434382 183218 446330 183454
rect 446566 183218 469826 183454
rect 434382 183134 469826 183218
rect 434382 182898 446330 183134
rect 446566 182898 469826 183134
rect 470382 183218 477050 183454
rect 477286 183218 505826 183454
rect 470382 183134 505826 183218
rect 470382 182898 477050 183134
rect 477286 182898 505826 183134
rect 506382 183218 507770 183454
rect 508006 183218 538490 183454
rect 538726 183218 541826 183454
rect 506382 183134 541826 183218
rect 506382 182898 507770 183134
rect 508006 182898 538490 183134
rect 538726 182898 541826 183134
rect 542382 183218 569210 183454
rect 569446 183218 577826 183454
rect 542382 183134 577826 183218
rect 542382 182898 569210 183134
rect 569446 182898 577826 183134
rect 578382 182898 585342 183454
rect 585898 182898 592650 183454
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 172938 -8694 173494
rect -8138 172938 27866 173494
rect 28422 172938 63866 173494
rect 64422 172938 99866 173494
rect 100422 172938 135866 173494
rect 136422 172938 171866 173494
rect 172422 172938 207866 173494
rect 208422 172938 243866 173494
rect 244422 172938 279866 173494
rect 280422 172938 315866 173494
rect 316422 172938 351866 173494
rect 352422 172938 387866 173494
rect 388422 172938 423866 173494
rect 424422 172938 459866 173494
rect 460422 172938 495866 173494
rect 496422 172938 531866 173494
rect 532422 172938 567866 173494
rect 568422 172938 592062 173494
rect 592618 172938 592650 173494
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169218 -7734 169774
rect -7178 169218 24146 169774
rect 24702 169218 60146 169774
rect 60702 169218 96146 169774
rect 96702 169218 132146 169774
rect 132702 169218 168146 169774
rect 168702 169218 204146 169774
rect 204702 169218 240146 169774
rect 240702 169218 276146 169774
rect 276702 169218 312146 169774
rect 312702 169218 348146 169774
rect 348702 169218 384146 169774
rect 384702 169218 420146 169774
rect 420702 169218 456146 169774
rect 456702 169218 528146 169774
rect 528702 169218 564146 169774
rect 564702 169218 591102 169774
rect 591658 169218 592650 169774
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165498 -6774 166054
rect -6218 165498 20426 166054
rect 20982 165498 56426 166054
rect 56982 165498 128426 166054
rect 128982 165498 164426 166054
rect 164982 165498 236426 166054
rect 236982 165498 272426 166054
rect 272982 165498 344426 166054
rect 344982 165498 380426 166054
rect 380982 165498 416426 166054
rect 416982 165498 452426 166054
rect 452982 165498 488426 166054
rect 488982 165498 524426 166054
rect 524982 165498 560426 166054
rect 560982 165498 590142 166054
rect 590698 165498 592650 166054
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 161778 -5814 162334
rect -5258 161778 16706 162334
rect 17262 161778 52706 162334
rect 53262 161778 88706 162334
rect 89262 161778 124706 162334
rect 125262 161778 160706 162334
rect 161262 161778 196706 162334
rect 197262 161778 232706 162334
rect 233262 161778 268706 162334
rect 269262 161778 304706 162334
rect 305262 161778 340706 162334
rect 341262 161778 376706 162334
rect 377262 161778 412706 162334
rect 413262 161778 448706 162334
rect 449262 161778 484706 162334
rect 485262 161778 520706 162334
rect 521262 161778 556706 162334
rect 557262 161778 589182 162334
rect 589738 161778 592650 162334
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158058 -4854 158614
rect -4298 158058 12986 158614
rect 13542 158058 48986 158614
rect 49542 158058 84986 158614
rect 85542 158058 120986 158614
rect 121542 158058 156986 158614
rect 157542 158058 192986 158614
rect 193542 158058 228986 158614
rect 229542 158058 264986 158614
rect 265542 158058 300986 158614
rect 301542 158058 336986 158614
rect 337542 158058 372986 158614
rect 373542 158058 408986 158614
rect 409542 158058 444986 158614
rect 445542 158058 480986 158614
rect 481542 158058 516986 158614
rect 517542 158058 552986 158614
rect 553542 158058 588222 158614
rect 588778 158058 592650 158614
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154338 -3894 154894
rect -3338 154338 9266 154894
rect 9822 154338 45266 154894
rect 45822 154338 81266 154894
rect 81822 154338 117266 154894
rect 117822 154338 153266 154894
rect 153822 154338 189266 154894
rect 189822 154338 225266 154894
rect 225822 154338 261266 154894
rect 261822 154338 297266 154894
rect 297822 154338 333266 154894
rect 333822 154338 405266 154894
rect 405822 154338 441266 154894
rect 441822 154338 513266 154894
rect 513822 154338 549266 154894
rect 549822 154338 587262 154894
rect 587818 154338 592650 154894
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150618 -2934 151174
rect -2378 150618 5546 151174
rect 6102 150938 31610 151174
rect 31846 150938 41546 151174
rect 6102 150854 41546 150938
rect 6102 150618 31610 150854
rect 31846 150618 41546 150854
rect 42102 150938 62330 151174
rect 62566 150938 93050 151174
rect 93286 150938 113546 151174
rect 42102 150854 113546 150938
rect 42102 150618 62330 150854
rect 62566 150618 93050 150854
rect 93286 150618 113546 150854
rect 114102 150938 123770 151174
rect 124006 150938 149546 151174
rect 114102 150854 149546 150938
rect 114102 150618 123770 150854
rect 124006 150618 149546 150854
rect 150102 150938 154490 151174
rect 154726 150938 185210 151174
rect 185446 150938 215930 151174
rect 216166 150938 221546 151174
rect 150102 150854 221546 150938
rect 150102 150618 154490 150854
rect 154726 150618 185210 150854
rect 185446 150618 215930 150854
rect 216166 150618 221546 150854
rect 222102 150938 246650 151174
rect 246886 150938 257546 151174
rect 222102 150854 257546 150938
rect 222102 150618 246650 150854
rect 246886 150618 257546 150854
rect 258102 150938 277370 151174
rect 277606 150938 293546 151174
rect 258102 150854 293546 150938
rect 258102 150618 277370 150854
rect 277606 150618 293546 150854
rect 294102 150938 308090 151174
rect 308326 150938 329546 151174
rect 294102 150854 329546 150938
rect 294102 150618 308090 150854
rect 308326 150618 329546 150854
rect 330102 150938 338810 151174
rect 339046 150938 365546 151174
rect 330102 150854 365546 150938
rect 330102 150618 338810 150854
rect 339046 150618 365546 150854
rect 366102 150938 369530 151174
rect 369766 150938 400250 151174
rect 400486 150938 401546 151174
rect 366102 150854 401546 150938
rect 366102 150618 369530 150854
rect 369766 150618 400250 150854
rect 400486 150618 401546 150854
rect 402102 150938 430970 151174
rect 431206 150938 437546 151174
rect 402102 150854 437546 150938
rect 402102 150618 430970 150854
rect 431206 150618 437546 150854
rect 438102 150938 461690 151174
rect 461926 150938 473546 151174
rect 438102 150854 473546 150938
rect 438102 150618 461690 150854
rect 461926 150618 473546 150854
rect 474102 150938 492410 151174
rect 492646 150938 509546 151174
rect 474102 150854 509546 150938
rect 474102 150618 492410 150854
rect 492646 150618 509546 150854
rect 510102 150938 523130 151174
rect 523366 150938 545546 151174
rect 510102 150854 545546 150938
rect 510102 150618 523130 150854
rect 523366 150618 545546 150854
rect 546102 150938 553850 151174
rect 554086 150938 581546 151174
rect 546102 150854 581546 150938
rect 546102 150618 553850 150854
rect 554086 150618 581546 150854
rect 582102 150618 586302 151174
rect 586858 150618 592650 151174
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 146898 -1974 147454
rect -1418 146898 1826 147454
rect 2382 147218 16250 147454
rect 16486 147218 37826 147454
rect 2382 147134 37826 147218
rect 2382 146898 16250 147134
rect 16486 146898 37826 147134
rect 38382 147218 46970 147454
rect 47206 147218 73826 147454
rect 38382 147134 73826 147218
rect 38382 146898 46970 147134
rect 47206 146898 73826 147134
rect 74382 147218 77690 147454
rect 77926 147218 108410 147454
rect 108646 147218 109826 147454
rect 74382 147134 109826 147218
rect 74382 146898 77690 147134
rect 77926 146898 108410 147134
rect 108646 146898 109826 147134
rect 110382 147218 139130 147454
rect 139366 147218 145826 147454
rect 110382 147134 145826 147218
rect 110382 146898 139130 147134
rect 139366 146898 145826 147134
rect 146382 147218 169850 147454
rect 170086 147218 181826 147454
rect 146382 147134 181826 147218
rect 146382 146898 169850 147134
rect 170086 146898 181826 147134
rect 182382 147218 200570 147454
rect 200806 147218 217826 147454
rect 182382 147134 217826 147218
rect 182382 146898 200570 147134
rect 200806 146898 217826 147134
rect 218382 147218 231290 147454
rect 231526 147218 253826 147454
rect 218382 147134 253826 147218
rect 218382 146898 231290 147134
rect 231526 146898 253826 147134
rect 254382 147218 262010 147454
rect 262246 147218 289826 147454
rect 254382 147134 289826 147218
rect 254382 146898 262010 147134
rect 262246 146898 289826 147134
rect 290382 147218 292730 147454
rect 292966 147218 323450 147454
rect 323686 147218 325826 147454
rect 290382 147134 325826 147218
rect 290382 146898 292730 147134
rect 292966 146898 323450 147134
rect 323686 146898 325826 147134
rect 326382 147218 354170 147454
rect 354406 147218 361826 147454
rect 326382 147134 361826 147218
rect 326382 146898 354170 147134
rect 354406 146898 361826 147134
rect 362382 147218 384890 147454
rect 385126 147218 397826 147454
rect 362382 147134 397826 147218
rect 362382 146898 384890 147134
rect 385126 146898 397826 147134
rect 398382 147218 415610 147454
rect 415846 147218 433826 147454
rect 398382 147134 433826 147218
rect 398382 146898 415610 147134
rect 415846 146898 433826 147134
rect 434382 147218 446330 147454
rect 446566 147218 469826 147454
rect 434382 147134 469826 147218
rect 434382 146898 446330 147134
rect 446566 146898 469826 147134
rect 470382 147218 477050 147454
rect 477286 147218 505826 147454
rect 470382 147134 505826 147218
rect 470382 146898 477050 147134
rect 477286 146898 505826 147134
rect 506382 147218 507770 147454
rect 508006 147218 538490 147454
rect 538726 147218 541826 147454
rect 506382 147134 541826 147218
rect 506382 146898 507770 147134
rect 508006 146898 538490 147134
rect 538726 146898 541826 147134
rect 542382 147218 569210 147454
rect 569446 147218 577826 147454
rect 542382 147134 577826 147218
rect 542382 146898 569210 147134
rect 569446 146898 577826 147134
rect 578382 146898 585342 147454
rect 585898 146898 592650 147454
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 136938 -8694 137494
rect -8138 136938 27866 137494
rect 28422 136938 63866 137494
rect 64422 136938 99866 137494
rect 100422 136938 135866 137494
rect 136422 136938 171866 137494
rect 172422 136938 207866 137494
rect 208422 136938 243866 137494
rect 244422 136938 279866 137494
rect 280422 136938 315866 137494
rect 316422 136938 351866 137494
rect 352422 136938 387866 137494
rect 388422 136938 423866 137494
rect 424422 136938 459866 137494
rect 460422 136938 495866 137494
rect 496422 136938 531866 137494
rect 532422 136938 567866 137494
rect 568422 136938 592062 137494
rect 592618 136938 592650 137494
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133218 -7734 133774
rect -7178 133218 24146 133774
rect 24702 133218 60146 133774
rect 60702 133218 96146 133774
rect 96702 133218 132146 133774
rect 132702 133218 168146 133774
rect 168702 133218 204146 133774
rect 204702 133218 240146 133774
rect 240702 133218 276146 133774
rect 276702 133218 312146 133774
rect 312702 133218 348146 133774
rect 348702 133218 384146 133774
rect 384702 133218 420146 133774
rect 420702 133218 456146 133774
rect 456702 133218 528146 133774
rect 528702 133218 564146 133774
rect 564702 133218 591102 133774
rect 591658 133218 592650 133774
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129498 -6774 130054
rect -6218 129498 20426 130054
rect 20982 129498 56426 130054
rect 56982 129498 128426 130054
rect 128982 129498 164426 130054
rect 164982 129498 236426 130054
rect 236982 129498 272426 130054
rect 272982 129498 344426 130054
rect 344982 129498 380426 130054
rect 380982 129498 416426 130054
rect 416982 129498 452426 130054
rect 452982 129498 488426 130054
rect 488982 129498 524426 130054
rect 524982 129498 560426 130054
rect 560982 129498 590142 130054
rect 590698 129498 592650 130054
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 125778 -5814 126334
rect -5258 125778 16706 126334
rect 17262 125778 52706 126334
rect 53262 125778 88706 126334
rect 89262 125778 124706 126334
rect 125262 125778 160706 126334
rect 161262 125778 196706 126334
rect 197262 125778 232706 126334
rect 233262 125778 268706 126334
rect 269262 125778 304706 126334
rect 305262 125778 340706 126334
rect 341262 125778 376706 126334
rect 377262 125778 412706 126334
rect 413262 125778 448706 126334
rect 449262 125778 484706 126334
rect 485262 125778 520706 126334
rect 521262 125778 556706 126334
rect 557262 125778 589182 126334
rect 589738 125778 592650 126334
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122058 -4854 122614
rect -4298 122058 12986 122614
rect 13542 122058 48986 122614
rect 49542 122058 84986 122614
rect 85542 122058 120986 122614
rect 121542 122058 156986 122614
rect 157542 122058 192986 122614
rect 193542 122058 228986 122614
rect 229542 122058 264986 122614
rect 265542 122058 300986 122614
rect 301542 122058 336986 122614
rect 337542 122058 372986 122614
rect 373542 122058 408986 122614
rect 409542 122058 444986 122614
rect 445542 122058 480986 122614
rect 481542 122058 516986 122614
rect 517542 122058 552986 122614
rect 553542 122058 588222 122614
rect 588778 122058 592650 122614
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118338 -3894 118894
rect -3338 118338 9266 118894
rect 9822 118338 45266 118894
rect 45822 118338 81266 118894
rect 81822 118338 117266 118894
rect 117822 118338 153266 118894
rect 153822 118338 189266 118894
rect 189822 118338 225266 118894
rect 225822 118338 261266 118894
rect 261822 118338 297266 118894
rect 297822 118338 333266 118894
rect 333822 118338 405266 118894
rect 405822 118338 441266 118894
rect 441822 118338 513266 118894
rect 513822 118338 549266 118894
rect 549822 118338 587262 118894
rect 587818 118338 592650 118894
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114618 -2934 115174
rect -2378 114618 5546 115174
rect 6102 114938 31610 115174
rect 31846 114938 41546 115174
rect 6102 114854 41546 114938
rect 6102 114618 31610 114854
rect 31846 114618 41546 114854
rect 42102 114938 62330 115174
rect 62566 114938 93050 115174
rect 93286 114938 113546 115174
rect 42102 114854 113546 114938
rect 42102 114618 62330 114854
rect 62566 114618 93050 114854
rect 93286 114618 113546 114854
rect 114102 114938 123770 115174
rect 124006 114938 149546 115174
rect 114102 114854 149546 114938
rect 114102 114618 123770 114854
rect 124006 114618 149546 114854
rect 150102 114938 154490 115174
rect 154726 114938 185210 115174
rect 185446 114938 215930 115174
rect 216166 114938 221546 115174
rect 150102 114854 221546 114938
rect 150102 114618 154490 114854
rect 154726 114618 185210 114854
rect 185446 114618 215930 114854
rect 216166 114618 221546 114854
rect 222102 114938 246650 115174
rect 246886 114938 257546 115174
rect 222102 114854 257546 114938
rect 222102 114618 246650 114854
rect 246886 114618 257546 114854
rect 258102 114938 277370 115174
rect 277606 114938 293546 115174
rect 258102 114854 293546 114938
rect 258102 114618 277370 114854
rect 277606 114618 293546 114854
rect 294102 114938 308090 115174
rect 308326 114938 329546 115174
rect 294102 114854 329546 114938
rect 294102 114618 308090 114854
rect 308326 114618 329546 114854
rect 330102 114938 338810 115174
rect 339046 114938 365546 115174
rect 330102 114854 365546 114938
rect 330102 114618 338810 114854
rect 339046 114618 365546 114854
rect 366102 114938 369530 115174
rect 369766 114938 400250 115174
rect 400486 114938 401546 115174
rect 366102 114854 401546 114938
rect 366102 114618 369530 114854
rect 369766 114618 400250 114854
rect 400486 114618 401546 114854
rect 402102 114938 430970 115174
rect 431206 114938 437546 115174
rect 402102 114854 437546 114938
rect 402102 114618 430970 114854
rect 431206 114618 437546 114854
rect 438102 114938 461690 115174
rect 461926 114938 473546 115174
rect 438102 114854 473546 114938
rect 438102 114618 461690 114854
rect 461926 114618 473546 114854
rect 474102 114938 492410 115174
rect 492646 114938 509546 115174
rect 474102 114854 509546 114938
rect 474102 114618 492410 114854
rect 492646 114618 509546 114854
rect 510102 114938 523130 115174
rect 523366 114938 545546 115174
rect 510102 114854 545546 114938
rect 510102 114618 523130 114854
rect 523366 114618 545546 114854
rect 546102 114938 553850 115174
rect 554086 114938 581546 115174
rect 546102 114854 581546 114938
rect 546102 114618 553850 114854
rect 554086 114618 581546 114854
rect 582102 114618 586302 115174
rect 586858 114618 592650 115174
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 110898 -1974 111454
rect -1418 110898 1826 111454
rect 2382 111218 16250 111454
rect 16486 111218 37826 111454
rect 2382 111134 37826 111218
rect 2382 110898 16250 111134
rect 16486 110898 37826 111134
rect 38382 111218 46970 111454
rect 47206 111218 73826 111454
rect 38382 111134 73826 111218
rect 38382 110898 46970 111134
rect 47206 110898 73826 111134
rect 74382 111218 77690 111454
rect 77926 111218 108410 111454
rect 108646 111218 109826 111454
rect 74382 111134 109826 111218
rect 74382 110898 77690 111134
rect 77926 110898 108410 111134
rect 108646 110898 109826 111134
rect 110382 111218 139130 111454
rect 139366 111218 145826 111454
rect 110382 111134 145826 111218
rect 110382 110898 139130 111134
rect 139366 110898 145826 111134
rect 146382 111218 169850 111454
rect 170086 111218 181826 111454
rect 146382 111134 181826 111218
rect 146382 110898 169850 111134
rect 170086 110898 181826 111134
rect 182382 111218 200570 111454
rect 200806 111218 217826 111454
rect 182382 111134 217826 111218
rect 182382 110898 200570 111134
rect 200806 110898 217826 111134
rect 218382 111218 231290 111454
rect 231526 111218 253826 111454
rect 218382 111134 253826 111218
rect 218382 110898 231290 111134
rect 231526 110898 253826 111134
rect 254382 111218 262010 111454
rect 262246 111218 289826 111454
rect 254382 111134 289826 111218
rect 254382 110898 262010 111134
rect 262246 110898 289826 111134
rect 290382 111218 292730 111454
rect 292966 111218 323450 111454
rect 323686 111218 325826 111454
rect 290382 111134 325826 111218
rect 290382 110898 292730 111134
rect 292966 110898 323450 111134
rect 323686 110898 325826 111134
rect 326382 111218 354170 111454
rect 354406 111218 361826 111454
rect 326382 111134 361826 111218
rect 326382 110898 354170 111134
rect 354406 110898 361826 111134
rect 362382 111218 384890 111454
rect 385126 111218 397826 111454
rect 362382 111134 397826 111218
rect 362382 110898 384890 111134
rect 385126 110898 397826 111134
rect 398382 111218 415610 111454
rect 415846 111218 433826 111454
rect 398382 111134 433826 111218
rect 398382 110898 415610 111134
rect 415846 110898 433826 111134
rect 434382 111218 446330 111454
rect 446566 111218 469826 111454
rect 434382 111134 469826 111218
rect 434382 110898 446330 111134
rect 446566 110898 469826 111134
rect 470382 111218 477050 111454
rect 477286 111218 505826 111454
rect 470382 111134 505826 111218
rect 470382 110898 477050 111134
rect 477286 110898 505826 111134
rect 506382 111218 507770 111454
rect 508006 111218 538490 111454
rect 538726 111218 541826 111454
rect 506382 111134 541826 111218
rect 506382 110898 507770 111134
rect 508006 110898 538490 111134
rect 538726 110898 541826 111134
rect 542382 111218 569210 111454
rect 569446 111218 577826 111454
rect 542382 111134 577826 111218
rect 542382 110898 569210 111134
rect 569446 110898 577826 111134
rect 578382 110898 585342 111454
rect 585898 110898 592650 111454
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 100938 -8694 101494
rect -8138 100938 27866 101494
rect 28422 100938 63866 101494
rect 64422 100938 99866 101494
rect 100422 100938 135866 101494
rect 136422 100938 171866 101494
rect 172422 100938 207866 101494
rect 208422 100938 243866 101494
rect 244422 100938 279866 101494
rect 280422 100938 315866 101494
rect 316422 100938 351866 101494
rect 352422 100938 387866 101494
rect 388422 100938 423866 101494
rect 424422 100938 459866 101494
rect 460422 100938 495866 101494
rect 496422 100938 531866 101494
rect 532422 100938 567866 101494
rect 568422 100938 592062 101494
rect 592618 100938 592650 101494
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97218 -7734 97774
rect -7178 97218 24146 97774
rect 24702 97218 60146 97774
rect 60702 97218 96146 97774
rect 96702 97218 132146 97774
rect 132702 97218 168146 97774
rect 168702 97218 204146 97774
rect 204702 97218 240146 97774
rect 240702 97218 276146 97774
rect 276702 97218 312146 97774
rect 312702 97218 348146 97774
rect 348702 97218 384146 97774
rect 384702 97218 420146 97774
rect 420702 97218 456146 97774
rect 456702 97218 528146 97774
rect 528702 97218 564146 97774
rect 564702 97218 591102 97774
rect 591658 97218 592650 97774
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93498 -6774 94054
rect -6218 93498 20426 94054
rect 20982 93498 56426 94054
rect 56982 93498 128426 94054
rect 128982 93498 164426 94054
rect 164982 93498 236426 94054
rect 236982 93498 272426 94054
rect 272982 93498 344426 94054
rect 344982 93498 380426 94054
rect 380982 93498 416426 94054
rect 416982 93498 452426 94054
rect 452982 93498 488426 94054
rect 488982 93498 524426 94054
rect 524982 93498 560426 94054
rect 560982 93498 590142 94054
rect 590698 93498 592650 94054
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 89778 -5814 90334
rect -5258 89778 16706 90334
rect 17262 89778 52706 90334
rect 53262 89778 88706 90334
rect 89262 89778 124706 90334
rect 125262 89778 160706 90334
rect 161262 89778 196706 90334
rect 197262 89778 232706 90334
rect 233262 89778 268706 90334
rect 269262 89778 304706 90334
rect 305262 89778 340706 90334
rect 341262 89778 376706 90334
rect 377262 89778 412706 90334
rect 413262 89778 448706 90334
rect 449262 89778 484706 90334
rect 485262 89778 520706 90334
rect 521262 89778 556706 90334
rect 557262 89778 589182 90334
rect 589738 89778 592650 90334
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86058 -4854 86614
rect -4298 86058 12986 86614
rect 13542 86058 48986 86614
rect 49542 86058 84986 86614
rect 85542 86058 120986 86614
rect 121542 86058 156986 86614
rect 157542 86058 192986 86614
rect 193542 86058 228986 86614
rect 229542 86058 264986 86614
rect 265542 86058 300986 86614
rect 301542 86058 336986 86614
rect 337542 86058 372986 86614
rect 373542 86058 408986 86614
rect 409542 86058 444986 86614
rect 445542 86058 480986 86614
rect 481542 86058 516986 86614
rect 517542 86058 552986 86614
rect 553542 86058 588222 86614
rect 588778 86058 592650 86614
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82338 -3894 82894
rect -3338 82338 9266 82894
rect 9822 82338 45266 82894
rect 45822 82338 81266 82894
rect 81822 82338 117266 82894
rect 117822 82338 153266 82894
rect 153822 82338 189266 82894
rect 189822 82338 225266 82894
rect 225822 82338 261266 82894
rect 261822 82338 297266 82894
rect 297822 82338 333266 82894
rect 333822 82338 405266 82894
rect 405822 82338 441266 82894
rect 441822 82338 513266 82894
rect 513822 82338 549266 82894
rect 549822 82338 587262 82894
rect 587818 82338 592650 82894
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78618 -2934 79174
rect -2378 78618 5546 79174
rect 6102 78938 31610 79174
rect 31846 78938 41546 79174
rect 6102 78854 41546 78938
rect 6102 78618 31610 78854
rect 31846 78618 41546 78854
rect 42102 78938 62330 79174
rect 62566 78938 93050 79174
rect 93286 78938 113546 79174
rect 42102 78854 113546 78938
rect 42102 78618 62330 78854
rect 62566 78618 93050 78854
rect 93286 78618 113546 78854
rect 114102 78938 123770 79174
rect 124006 78938 149546 79174
rect 114102 78854 149546 78938
rect 114102 78618 123770 78854
rect 124006 78618 149546 78854
rect 150102 78938 154490 79174
rect 154726 78938 185210 79174
rect 185446 78938 215930 79174
rect 216166 78938 221546 79174
rect 150102 78854 221546 78938
rect 150102 78618 154490 78854
rect 154726 78618 185210 78854
rect 185446 78618 215930 78854
rect 216166 78618 221546 78854
rect 222102 78938 246650 79174
rect 246886 78938 257546 79174
rect 222102 78854 257546 78938
rect 222102 78618 246650 78854
rect 246886 78618 257546 78854
rect 258102 78938 277370 79174
rect 277606 78938 293546 79174
rect 258102 78854 293546 78938
rect 258102 78618 277370 78854
rect 277606 78618 293546 78854
rect 294102 78938 308090 79174
rect 308326 78938 329546 79174
rect 294102 78854 329546 78938
rect 294102 78618 308090 78854
rect 308326 78618 329546 78854
rect 330102 78938 338810 79174
rect 339046 78938 365546 79174
rect 330102 78854 365546 78938
rect 330102 78618 338810 78854
rect 339046 78618 365546 78854
rect 366102 78938 369530 79174
rect 369766 78938 400250 79174
rect 400486 78938 401546 79174
rect 366102 78854 401546 78938
rect 366102 78618 369530 78854
rect 369766 78618 400250 78854
rect 400486 78618 401546 78854
rect 402102 78938 430970 79174
rect 431206 78938 437546 79174
rect 402102 78854 437546 78938
rect 402102 78618 430970 78854
rect 431206 78618 437546 78854
rect 438102 78938 461690 79174
rect 461926 78938 473546 79174
rect 438102 78854 473546 78938
rect 438102 78618 461690 78854
rect 461926 78618 473546 78854
rect 474102 78938 492410 79174
rect 492646 78938 509546 79174
rect 474102 78854 509546 78938
rect 474102 78618 492410 78854
rect 492646 78618 509546 78854
rect 510102 78938 523130 79174
rect 523366 78938 545546 79174
rect 510102 78854 545546 78938
rect 510102 78618 523130 78854
rect 523366 78618 545546 78854
rect 546102 78938 553850 79174
rect 554086 78938 581546 79174
rect 546102 78854 581546 78938
rect 546102 78618 553850 78854
rect 554086 78618 581546 78854
rect 582102 78618 586302 79174
rect 586858 78618 592650 79174
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 74898 -1974 75454
rect -1418 74898 1826 75454
rect 2382 75218 16250 75454
rect 16486 75218 37826 75454
rect 2382 75134 37826 75218
rect 2382 74898 16250 75134
rect 16486 74898 37826 75134
rect 38382 75218 46970 75454
rect 47206 75218 73826 75454
rect 38382 75134 73826 75218
rect 38382 74898 46970 75134
rect 47206 74898 73826 75134
rect 74382 75218 77690 75454
rect 77926 75218 108410 75454
rect 108646 75218 109826 75454
rect 74382 75134 109826 75218
rect 74382 74898 77690 75134
rect 77926 74898 108410 75134
rect 108646 74898 109826 75134
rect 110382 75218 139130 75454
rect 139366 75218 145826 75454
rect 110382 75134 145826 75218
rect 110382 74898 139130 75134
rect 139366 74898 145826 75134
rect 146382 75218 169850 75454
rect 170086 75218 181826 75454
rect 146382 75134 181826 75218
rect 146382 74898 169850 75134
rect 170086 74898 181826 75134
rect 182382 75218 200570 75454
rect 200806 75218 217826 75454
rect 182382 75134 217826 75218
rect 182382 74898 200570 75134
rect 200806 74898 217826 75134
rect 218382 75218 231290 75454
rect 231526 75218 253826 75454
rect 218382 75134 253826 75218
rect 218382 74898 231290 75134
rect 231526 74898 253826 75134
rect 254382 75218 262010 75454
rect 262246 75218 289826 75454
rect 254382 75134 289826 75218
rect 254382 74898 262010 75134
rect 262246 74898 289826 75134
rect 290382 75218 292730 75454
rect 292966 75218 323450 75454
rect 323686 75218 325826 75454
rect 290382 75134 325826 75218
rect 290382 74898 292730 75134
rect 292966 74898 323450 75134
rect 323686 74898 325826 75134
rect 326382 75218 354170 75454
rect 354406 75218 361826 75454
rect 326382 75134 361826 75218
rect 326382 74898 354170 75134
rect 354406 74898 361826 75134
rect 362382 75218 384890 75454
rect 385126 75218 397826 75454
rect 362382 75134 397826 75218
rect 362382 74898 384890 75134
rect 385126 74898 397826 75134
rect 398382 75218 415610 75454
rect 415846 75218 433826 75454
rect 398382 75134 433826 75218
rect 398382 74898 415610 75134
rect 415846 74898 433826 75134
rect 434382 75218 446330 75454
rect 446566 75218 469826 75454
rect 434382 75134 469826 75218
rect 434382 74898 446330 75134
rect 446566 74898 469826 75134
rect 470382 75218 477050 75454
rect 477286 75218 505826 75454
rect 470382 75134 505826 75218
rect 470382 74898 477050 75134
rect 477286 74898 505826 75134
rect 506382 75218 507770 75454
rect 508006 75218 538490 75454
rect 538726 75218 541826 75454
rect 506382 75134 541826 75218
rect 506382 74898 507770 75134
rect 508006 74898 538490 75134
rect 538726 74898 541826 75134
rect 542382 75218 569210 75454
rect 569446 75218 577826 75454
rect 542382 75134 577826 75218
rect 542382 74898 569210 75134
rect 569446 74898 577826 75134
rect 578382 74898 585342 75454
rect 585898 74898 592650 75454
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 64938 -8694 65494
rect -8138 64938 27866 65494
rect 28422 64938 63866 65494
rect 64422 64938 99866 65494
rect 100422 64938 135866 65494
rect 136422 64938 171866 65494
rect 172422 64938 207866 65494
rect 208422 64938 243866 65494
rect 244422 64938 279866 65494
rect 280422 64938 315866 65494
rect 316422 64938 351866 65494
rect 352422 64938 387866 65494
rect 388422 64938 423866 65494
rect 424422 64938 459866 65494
rect 460422 64938 495866 65494
rect 496422 64938 531866 65494
rect 532422 64938 567866 65494
rect 568422 64938 592062 65494
rect 592618 64938 592650 65494
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61218 -7734 61774
rect -7178 61218 24146 61774
rect 24702 61218 60146 61774
rect 60702 61218 96146 61774
rect 96702 61218 132146 61774
rect 132702 61218 168146 61774
rect 168702 61218 204146 61774
rect 204702 61218 240146 61774
rect 240702 61218 276146 61774
rect 276702 61218 312146 61774
rect 312702 61218 348146 61774
rect 348702 61218 384146 61774
rect 384702 61218 420146 61774
rect 420702 61218 456146 61774
rect 456702 61218 528146 61774
rect 528702 61218 564146 61774
rect 564702 61218 591102 61774
rect 591658 61218 592650 61774
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57498 -6774 58054
rect -6218 57498 20426 58054
rect 20982 57498 56426 58054
rect 56982 57498 128426 58054
rect 128982 57498 164426 58054
rect 164982 57498 236426 58054
rect 236982 57498 272426 58054
rect 272982 57498 344426 58054
rect 344982 57498 380426 58054
rect 380982 57498 416426 58054
rect 416982 57498 452426 58054
rect 452982 57498 488426 58054
rect 488982 57498 524426 58054
rect 524982 57498 560426 58054
rect 560982 57498 590142 58054
rect 590698 57498 592650 58054
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 53778 -5814 54334
rect -5258 53778 16706 54334
rect 17262 53778 52706 54334
rect 53262 53778 88706 54334
rect 89262 53778 124706 54334
rect 125262 53778 160706 54334
rect 161262 53778 196706 54334
rect 197262 53778 232706 54334
rect 233262 53778 268706 54334
rect 269262 53778 304706 54334
rect 305262 53778 340706 54334
rect 341262 53778 376706 54334
rect 377262 53778 412706 54334
rect 413262 53778 448706 54334
rect 449262 53778 484706 54334
rect 485262 53778 520706 54334
rect 521262 53778 556706 54334
rect 557262 53778 589182 54334
rect 589738 53778 592650 54334
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50058 -4854 50614
rect -4298 50058 12986 50614
rect 13542 50058 48986 50614
rect 49542 50058 84986 50614
rect 85542 50058 120986 50614
rect 121542 50058 156986 50614
rect 157542 50058 192986 50614
rect 193542 50058 228986 50614
rect 229542 50058 264986 50614
rect 265542 50058 300986 50614
rect 301542 50058 336986 50614
rect 337542 50058 372986 50614
rect 373542 50058 408986 50614
rect 409542 50058 444986 50614
rect 445542 50058 480986 50614
rect 481542 50058 516986 50614
rect 517542 50058 552986 50614
rect 553542 50058 588222 50614
rect 588778 50058 592650 50614
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46338 -3894 46894
rect -3338 46338 9266 46894
rect 9822 46338 45266 46894
rect 45822 46338 81266 46894
rect 81822 46338 117266 46894
rect 117822 46338 153266 46894
rect 153822 46338 189266 46894
rect 189822 46338 225266 46894
rect 225822 46338 261266 46894
rect 261822 46338 297266 46894
rect 297822 46338 333266 46894
rect 333822 46338 405266 46894
rect 405822 46338 441266 46894
rect 441822 46338 513266 46894
rect 513822 46338 549266 46894
rect 549822 46338 587262 46894
rect 587818 46338 592650 46894
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42618 -2934 43174
rect -2378 42618 5546 43174
rect 6102 42938 31610 43174
rect 31846 42938 41546 43174
rect 6102 42854 41546 42938
rect 6102 42618 31610 42854
rect 31846 42618 41546 42854
rect 42102 42938 62330 43174
rect 62566 42938 93050 43174
rect 93286 42938 113546 43174
rect 42102 42854 113546 42938
rect 42102 42618 62330 42854
rect 62566 42618 93050 42854
rect 93286 42618 113546 42854
rect 114102 42938 123770 43174
rect 124006 42938 149546 43174
rect 114102 42854 149546 42938
rect 114102 42618 123770 42854
rect 124006 42618 149546 42854
rect 150102 42938 154490 43174
rect 154726 42938 185210 43174
rect 185446 42938 215930 43174
rect 216166 42938 221546 43174
rect 150102 42854 221546 42938
rect 150102 42618 154490 42854
rect 154726 42618 185210 42854
rect 185446 42618 215930 42854
rect 216166 42618 221546 42854
rect 222102 42938 246650 43174
rect 246886 42938 257546 43174
rect 222102 42854 257546 42938
rect 222102 42618 246650 42854
rect 246886 42618 257546 42854
rect 258102 42938 277370 43174
rect 277606 42938 293546 43174
rect 258102 42854 293546 42938
rect 258102 42618 277370 42854
rect 277606 42618 293546 42854
rect 294102 42938 308090 43174
rect 308326 42938 329546 43174
rect 294102 42854 329546 42938
rect 294102 42618 308090 42854
rect 308326 42618 329546 42854
rect 330102 42938 338810 43174
rect 339046 42938 365546 43174
rect 330102 42854 365546 42938
rect 330102 42618 338810 42854
rect 339046 42618 365546 42854
rect 366102 42938 369530 43174
rect 369766 42938 400250 43174
rect 400486 42938 401546 43174
rect 366102 42854 401546 42938
rect 366102 42618 369530 42854
rect 369766 42618 400250 42854
rect 400486 42618 401546 42854
rect 402102 42938 430970 43174
rect 431206 42938 437546 43174
rect 402102 42854 437546 42938
rect 402102 42618 430970 42854
rect 431206 42618 437546 42854
rect 438102 42938 461690 43174
rect 461926 42938 473546 43174
rect 438102 42854 473546 42938
rect 438102 42618 461690 42854
rect 461926 42618 473546 42854
rect 474102 42938 492410 43174
rect 492646 42938 509546 43174
rect 474102 42854 509546 42938
rect 474102 42618 492410 42854
rect 492646 42618 509546 42854
rect 510102 42938 523130 43174
rect 523366 42938 545546 43174
rect 510102 42854 545546 42938
rect 510102 42618 523130 42854
rect 523366 42618 545546 42854
rect 546102 42938 553850 43174
rect 554086 42938 581546 43174
rect 546102 42854 581546 42938
rect 546102 42618 553850 42854
rect 554086 42618 581546 42854
rect 582102 42618 586302 43174
rect 586858 42618 592650 43174
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 38898 -1974 39454
rect -1418 38898 1826 39454
rect 2382 39218 16250 39454
rect 16486 39218 37826 39454
rect 2382 39134 37826 39218
rect 2382 38898 16250 39134
rect 16486 38898 37826 39134
rect 38382 39218 46970 39454
rect 47206 39218 73826 39454
rect 38382 39134 73826 39218
rect 38382 38898 46970 39134
rect 47206 38898 73826 39134
rect 74382 39218 77690 39454
rect 77926 39218 108410 39454
rect 108646 39218 109826 39454
rect 74382 39134 109826 39218
rect 74382 38898 77690 39134
rect 77926 38898 108410 39134
rect 108646 38898 109826 39134
rect 110382 39218 139130 39454
rect 139366 39218 145826 39454
rect 110382 39134 145826 39218
rect 110382 38898 139130 39134
rect 139366 38898 145826 39134
rect 146382 39218 169850 39454
rect 170086 39218 181826 39454
rect 146382 39134 181826 39218
rect 146382 38898 169850 39134
rect 170086 38898 181826 39134
rect 182382 39218 200570 39454
rect 200806 39218 217826 39454
rect 182382 39134 217826 39218
rect 182382 38898 200570 39134
rect 200806 38898 217826 39134
rect 218382 39218 231290 39454
rect 231526 39218 253826 39454
rect 218382 39134 253826 39218
rect 218382 38898 231290 39134
rect 231526 38898 253826 39134
rect 254382 39218 262010 39454
rect 262246 39218 289826 39454
rect 254382 39134 289826 39218
rect 254382 38898 262010 39134
rect 262246 38898 289826 39134
rect 290382 39218 292730 39454
rect 292966 39218 323450 39454
rect 323686 39218 325826 39454
rect 290382 39134 325826 39218
rect 290382 38898 292730 39134
rect 292966 38898 323450 39134
rect 323686 38898 325826 39134
rect 326382 39218 354170 39454
rect 354406 39218 361826 39454
rect 326382 39134 361826 39218
rect 326382 38898 354170 39134
rect 354406 38898 361826 39134
rect 362382 39218 384890 39454
rect 385126 39218 397826 39454
rect 362382 39134 397826 39218
rect 362382 38898 384890 39134
rect 385126 38898 397826 39134
rect 398382 39218 415610 39454
rect 415846 39218 433826 39454
rect 398382 39134 433826 39218
rect 398382 38898 415610 39134
rect 415846 38898 433826 39134
rect 434382 39218 446330 39454
rect 446566 39218 469826 39454
rect 434382 39134 469826 39218
rect 434382 38898 446330 39134
rect 446566 38898 469826 39134
rect 470382 39218 477050 39454
rect 477286 39218 505826 39454
rect 470382 39134 505826 39218
rect 470382 38898 477050 39134
rect 477286 38898 505826 39134
rect 506382 39218 507770 39454
rect 508006 39218 538490 39454
rect 538726 39218 541826 39454
rect 506382 39134 541826 39218
rect 506382 38898 507770 39134
rect 508006 38898 538490 39134
rect 538726 38898 541826 39134
rect 542382 39218 569210 39454
rect 569446 39218 577826 39454
rect 542382 39134 577826 39218
rect 542382 38898 569210 39134
rect 569446 38898 577826 39134
rect 578382 38898 585342 39454
rect 585898 38898 592650 39454
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 28938 -8694 29494
rect -8138 28938 27866 29494
rect 28422 28938 63866 29494
rect 64422 28938 99866 29494
rect 100422 28938 135866 29494
rect 136422 28938 171866 29494
rect 172422 28938 207866 29494
rect 208422 28938 243866 29494
rect 244422 28938 279866 29494
rect 280422 28938 315866 29494
rect 316422 28938 351866 29494
rect 352422 28938 387866 29494
rect 388422 28938 423866 29494
rect 424422 28938 459866 29494
rect 460422 28938 495866 29494
rect 496422 28938 531866 29494
rect 532422 28938 567866 29494
rect 568422 28938 592062 29494
rect 592618 28938 592650 29494
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25218 -7734 25774
rect -7178 25218 24146 25774
rect 24702 25218 60146 25774
rect 60702 25218 96146 25774
rect 96702 25218 132146 25774
rect 132702 25218 168146 25774
rect 168702 25218 204146 25774
rect 204702 25218 276146 25774
rect 276702 25218 312146 25774
rect 312702 25218 348146 25774
rect 348702 25218 384146 25774
rect 384702 25218 420146 25774
rect 420702 25218 456146 25774
rect 456702 25218 528146 25774
rect 528702 25218 564146 25774
rect 564702 25218 591102 25774
rect 591658 25218 592650 25774
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21498 -6774 22054
rect -6218 21498 20426 22054
rect 20982 21498 56426 22054
rect 56982 21498 128426 22054
rect 128982 21498 164426 22054
rect 164982 21498 236426 22054
rect 236982 21498 272426 22054
rect 272982 21498 344426 22054
rect 344982 21498 380426 22054
rect 380982 21498 416426 22054
rect 416982 21498 452426 22054
rect 452982 21498 488426 22054
rect 488982 21498 524426 22054
rect 524982 21498 560426 22054
rect 560982 21498 590142 22054
rect 590698 21498 592650 22054
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 17778 -5814 18334
rect -5258 17778 16706 18334
rect 17262 17778 52706 18334
rect 53262 17778 88706 18334
rect 89262 17778 124706 18334
rect 125262 17778 160706 18334
rect 161262 17778 196706 18334
rect 197262 17778 232706 18334
rect 233262 17778 268706 18334
rect 269262 17778 304706 18334
rect 305262 17778 340706 18334
rect 341262 17778 376706 18334
rect 377262 17778 412706 18334
rect 413262 17778 448706 18334
rect 449262 17778 484706 18334
rect 485262 17778 520706 18334
rect 521262 17778 556706 18334
rect 557262 17778 589182 18334
rect 589738 17778 592650 18334
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14058 -4854 14614
rect -4298 14058 12986 14614
rect 13542 14058 48986 14614
rect 49542 14058 84986 14614
rect 85542 14058 120986 14614
rect 121542 14058 156986 14614
rect 157542 14058 192986 14614
rect 193542 14058 228986 14614
rect 229542 14058 264986 14614
rect 265542 14058 300986 14614
rect 301542 14058 336986 14614
rect 337542 14058 372986 14614
rect 373542 14058 408986 14614
rect 409542 14058 444986 14614
rect 445542 14058 480986 14614
rect 481542 14058 516986 14614
rect 517542 14058 552986 14614
rect 553542 14058 588222 14614
rect 588778 14058 592650 14614
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10338 -3894 10894
rect -3338 10338 9266 10894
rect 9822 10338 45266 10894
rect 45822 10338 81266 10894
rect 81822 10338 117266 10894
rect 117822 10338 153266 10894
rect 153822 10338 189266 10894
rect 189822 10338 225266 10894
rect 225822 10338 261266 10894
rect 261822 10338 297266 10894
rect 297822 10338 333266 10894
rect 333822 10338 405266 10894
rect 405822 10338 441266 10894
rect 441822 10338 513266 10894
rect 513822 10338 549266 10894
rect 549822 10338 587262 10894
rect 587818 10338 592650 10894
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6618 -2934 7174
rect -2378 6618 5546 7174
rect 6102 6938 31610 7174
rect 31846 6938 41546 7174
rect 6102 6854 41546 6938
rect 6102 6618 31610 6854
rect 31846 6618 41546 6854
rect 42102 6938 62330 7174
rect 62566 6938 93050 7174
rect 93286 6938 113546 7174
rect 42102 6854 113546 6938
rect 42102 6618 62330 6854
rect 62566 6618 93050 6854
rect 93286 6618 113546 6854
rect 114102 6938 123770 7174
rect 124006 6938 149546 7174
rect 114102 6854 149546 6938
rect 114102 6618 123770 6854
rect 124006 6618 149546 6854
rect 150102 6938 154490 7174
rect 154726 6938 185210 7174
rect 185446 6938 215930 7174
rect 216166 6938 221546 7174
rect 150102 6854 221546 6938
rect 150102 6618 154490 6854
rect 154726 6618 185210 6854
rect 185446 6618 215930 6854
rect 216166 6618 221546 6854
rect 222102 6938 246650 7174
rect 246886 6938 277370 7174
rect 277606 6938 293546 7174
rect 222102 6854 293546 6938
rect 222102 6618 246650 6854
rect 246886 6618 277370 6854
rect 277606 6618 293546 6854
rect 294102 6938 308090 7174
rect 308326 6938 329546 7174
rect 294102 6854 329546 6938
rect 294102 6618 308090 6854
rect 308326 6618 329546 6854
rect 330102 6938 338810 7174
rect 339046 6938 365546 7174
rect 330102 6854 365546 6938
rect 330102 6618 338810 6854
rect 339046 6618 365546 6854
rect 366102 6938 369530 7174
rect 369766 6938 400250 7174
rect 400486 6938 401546 7174
rect 366102 6854 401546 6938
rect 366102 6618 369530 6854
rect 369766 6618 400250 6854
rect 400486 6618 401546 6854
rect 402102 6938 430970 7174
rect 431206 6938 437546 7174
rect 402102 6854 437546 6938
rect 402102 6618 430970 6854
rect 431206 6618 437546 6854
rect 438102 6938 461690 7174
rect 461926 6938 473546 7174
rect 438102 6854 473546 6938
rect 438102 6618 461690 6854
rect 461926 6618 473546 6854
rect 474102 6938 492410 7174
rect 492646 6938 509546 7174
rect 474102 6854 509546 6938
rect 474102 6618 492410 6854
rect 492646 6618 509546 6854
rect 510102 6938 523130 7174
rect 523366 6938 545546 7174
rect 510102 6854 545546 6938
rect 510102 6618 523130 6854
rect 523366 6618 545546 6854
rect 546102 6938 553850 7174
rect 554086 6938 581546 7174
rect 546102 6854 581546 6938
rect 546102 6618 553850 6854
rect 554086 6618 581546 6854
rect 582102 6618 586302 7174
rect 586858 6618 592650 7174
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 2898 -1974 3454
rect -1418 2898 1826 3454
rect 2382 2898 37826 3454
rect 38382 2898 73826 3454
rect 74382 2898 109826 3454
rect 110382 2898 145826 3454
rect 146382 2898 181826 3454
rect 182382 2898 217826 3454
rect 218382 2898 253826 3454
rect 254382 2898 289826 3454
rect 290382 2898 325826 3454
rect 326382 2898 361826 3454
rect 362382 2898 397826 3454
rect 398382 2898 433826 3454
rect 434382 2898 469826 3454
rect 470382 2898 505826 3454
rect 506382 2898 541826 3454
rect 542382 2898 577826 3454
rect 578382 2898 585342 3454
rect 585898 2898 592650 3454
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -902 -1974 -346
rect -1418 -902 1826 -346
rect 2382 -902 37826 -346
rect 38382 -902 73826 -346
rect 74382 -902 109826 -346
rect 110382 -902 145826 -346
rect 146382 -902 181826 -346
rect 182382 -902 217826 -346
rect 218382 -902 253826 -346
rect 254382 -902 289826 -346
rect 290382 -902 325826 -346
rect 326382 -902 361826 -346
rect 362382 -902 397826 -346
rect 398382 -902 433826 -346
rect 434382 -902 469826 -346
rect 470382 -902 505826 -346
rect 506382 -902 541826 -346
rect 542382 -902 577826 -346
rect 578382 -902 585342 -346
rect 585898 -902 585930 -346
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1862 -2934 -1306
rect -2378 -1862 5546 -1306
rect 6102 -1862 41546 -1306
rect 42102 -1862 113546 -1306
rect 114102 -1862 149546 -1306
rect 150102 -1862 221546 -1306
rect 222102 -1862 293546 -1306
rect 294102 -1862 329546 -1306
rect 330102 -1862 365546 -1306
rect 366102 -1862 401546 -1306
rect 402102 -1862 437546 -1306
rect 438102 -1862 473546 -1306
rect 474102 -1862 509546 -1306
rect 510102 -1862 545546 -1306
rect 546102 -1862 581546 -1306
rect 582102 -1862 586302 -1306
rect 586858 -1862 586890 -1306
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2822 -3894 -2266
rect -3338 -2822 9266 -2266
rect 9822 -2822 45266 -2266
rect 45822 -2822 81266 -2266
rect 81822 -2822 117266 -2266
rect 117822 -2822 153266 -2266
rect 153822 -2822 189266 -2266
rect 189822 -2822 225266 -2266
rect 225822 -2822 261266 -2266
rect 261822 -2822 297266 -2266
rect 297822 -2822 333266 -2266
rect 333822 -2822 405266 -2266
rect 405822 -2822 441266 -2266
rect 441822 -2822 513266 -2266
rect 513822 -2822 549266 -2266
rect 549822 -2822 587262 -2266
rect 587818 -2822 587850 -2266
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3782 -4854 -3226
rect -4298 -3782 12986 -3226
rect 13542 -3782 48986 -3226
rect 49542 -3782 84986 -3226
rect 85542 -3782 120986 -3226
rect 121542 -3782 156986 -3226
rect 157542 -3782 192986 -3226
rect 193542 -3782 228986 -3226
rect 229542 -3782 264986 -3226
rect 265542 -3782 300986 -3226
rect 301542 -3782 336986 -3226
rect 337542 -3782 372986 -3226
rect 373542 -3782 408986 -3226
rect 409542 -3782 444986 -3226
rect 445542 -3782 480986 -3226
rect 481542 -3782 516986 -3226
rect 517542 -3782 552986 -3226
rect 553542 -3782 588222 -3226
rect 588778 -3782 588810 -3226
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4742 -5814 -4186
rect -5258 -4742 16706 -4186
rect 17262 -4742 52706 -4186
rect 53262 -4742 88706 -4186
rect 89262 -4742 124706 -4186
rect 125262 -4742 160706 -4186
rect 161262 -4742 196706 -4186
rect 197262 -4742 232706 -4186
rect 233262 -4742 268706 -4186
rect 269262 -4742 304706 -4186
rect 305262 -4742 340706 -4186
rect 341262 -4742 376706 -4186
rect 377262 -4742 412706 -4186
rect 413262 -4742 448706 -4186
rect 449262 -4742 484706 -4186
rect 485262 -4742 520706 -4186
rect 521262 -4742 556706 -4186
rect 557262 -4742 589182 -4186
rect 589738 -4742 589770 -4186
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5702 -6774 -5146
rect -6218 -5702 20426 -5146
rect 20982 -5702 56426 -5146
rect 56982 -5702 128426 -5146
rect 128982 -5702 164426 -5146
rect 164982 -5702 236426 -5146
rect 236982 -5702 272426 -5146
rect 272982 -5702 344426 -5146
rect 344982 -5702 380426 -5146
rect 380982 -5702 416426 -5146
rect 416982 -5702 452426 -5146
rect 452982 -5702 488426 -5146
rect 488982 -5702 524426 -5146
rect 524982 -5702 560426 -5146
rect 560982 -5702 590142 -5146
rect 590698 -5702 590730 -5146
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6662 -7734 -6106
rect -7178 -6662 24146 -6106
rect 24702 -6662 60146 -6106
rect 60702 -6662 96146 -6106
rect 96702 -6662 132146 -6106
rect 132702 -6662 168146 -6106
rect 168702 -6662 204146 -6106
rect 204702 -6662 276146 -6106
rect 276702 -6662 312146 -6106
rect 312702 -6662 348146 -6106
rect 348702 -6662 384146 -6106
rect 384702 -6662 420146 -6106
rect 420702 -6662 456146 -6106
rect 456702 -6662 528146 -6106
rect 528702 -6662 564146 -6106
rect 564702 -6662 591102 -6106
rect 591658 -6662 591690 -6106
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7622 -8694 -7066
rect -8138 -7622 27866 -7066
rect 28422 -7622 63866 -7066
rect 64422 -7622 99866 -7066
rect 100422 -7622 135866 -7066
rect 136422 -7622 171866 -7066
rect 172422 -7622 207866 -7066
rect 208422 -7622 279866 -7066
rect 280422 -7622 315866 -7066
rect 316422 -7622 351866 -7066
rect 352422 -7622 387866 -7066
rect 388422 -7622 423866 -7066
rect 424422 -7622 459866 -7066
rect 460422 -7622 495866 -7066
rect 496422 -7622 531866 -7066
rect 532422 -7622 567866 -7066
rect 568422 -7622 592062 -7066
rect 592618 -7622 592650 -7066
rect -8726 -7654 592650 -7622
use user_proj_example  mprj
timestamp 0
transform 1 0 12000 0 1 3000
box 0 0 560000 349840
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 1200 0 0 0 analog_io[0]
port 1 nsew
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 560 90 0 0 analog_io[10]
port 2 nsew
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 560 90 0 0 analog_io[11]
port 3 nsew
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 560 90 0 0 analog_io[12]
port 4 nsew
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 560 90 0 0 analog_io[13]
port 5 nsew
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 560 90 0 0 analog_io[14]
port 6 nsew
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 560 90 0 0 analog_io[15]
port 7 nsew
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 560 90 0 0 analog_io[16]
port 8 nsew
flabel metal3 s -960 697220 480 697460 0 FreeSans 1200 0 0 0 analog_io[17]
port 9 nsew
flabel metal3 s -960 644996 480 645236 0 FreeSans 1200 0 0 0 analog_io[18]
port 10 nsew
flabel metal3 s -960 592908 480 593148 0 FreeSans 1200 0 0 0 analog_io[19]
port 11 nsew
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 1200 0 0 0 analog_io[1]
port 12 nsew
flabel metal3 s -960 540684 480 540924 0 FreeSans 1200 0 0 0 analog_io[20]
port 13 nsew
flabel metal3 s -960 488596 480 488836 0 FreeSans 1200 0 0 0 analog_io[21]
port 14 nsew
flabel metal3 s -960 436508 480 436748 0 FreeSans 1200 0 0 0 analog_io[22]
port 15 nsew
flabel metal3 s -960 384284 480 384524 0 FreeSans 1200 0 0 0 analog_io[23]
port 16 nsew
flabel metal3 s -960 332196 480 332436 0 FreeSans 1200 0 0 0 analog_io[24]
port 17 nsew
flabel metal3 s -960 279972 480 280212 0 FreeSans 1200 0 0 0 analog_io[25]
port 18 nsew
flabel metal3 s -960 227884 480 228124 0 FreeSans 1200 0 0 0 analog_io[26]
port 19 nsew
flabel metal3 s -960 175796 480 176036 0 FreeSans 1200 0 0 0 analog_io[27]
port 20 nsew
flabel metal3 s -960 123572 480 123812 0 FreeSans 1200 0 0 0 analog_io[28]
port 21 nsew
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 1200 0 0 0 analog_io[2]
port 22 nsew
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 1200 0 0 0 analog_io[3]
port 23 nsew
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 1200 0 0 0 analog_io[4]
port 24 nsew
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 1200 0 0 0 analog_io[5]
port 25 nsew
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 1200 0 0 0 analog_io[6]
port 26 nsew
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 1200 0 0 0 analog_io[7]
port 27 nsew
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 560 90 0 0 analog_io[8]
port 28 nsew
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 560 90 0 0 analog_io[9]
port 29 nsew
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 1200 0 0 0 io_in[0]
port 30 nsew
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 1200 0 0 0 io_in[10]
port 31 nsew
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 1200 0 0 0 io_in[11]
port 32 nsew
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 1200 0 0 0 io_in[12]
port 33 nsew
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 1200 0 0 0 io_in[13]
port 34 nsew
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 1200 0 0 0 io_in[14]
port 35 nsew
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 560 90 0 0 io_in[15]
port 36 nsew
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 560 90 0 0 io_in[16]
port 37 nsew
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 560 90 0 0 io_in[17]
port 38 nsew
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 560 90 0 0 io_in[18]
port 39 nsew
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 560 90 0 0 io_in[19]
port 40 nsew
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 1200 0 0 0 io_in[1]
port 41 nsew
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 560 90 0 0 io_in[20]
port 42 nsew
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 560 90 0 0 io_in[21]
port 43 nsew
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 560 90 0 0 io_in[22]
port 44 nsew
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 560 90 0 0 io_in[23]
port 45 nsew
flabel metal3 s -960 684164 480 684404 0 FreeSans 1200 0 0 0 io_in[24]
port 46 nsew
flabel metal3 s -960 631940 480 632180 0 FreeSans 1200 0 0 0 io_in[25]
port 47 nsew
flabel metal3 s -960 579852 480 580092 0 FreeSans 1200 0 0 0 io_in[26]
port 48 nsew
flabel metal3 s -960 527764 480 528004 0 FreeSans 1200 0 0 0 io_in[27]
port 49 nsew
flabel metal3 s -960 475540 480 475780 0 FreeSans 1200 0 0 0 io_in[28]
port 50 nsew
flabel metal3 s -960 423452 480 423692 0 FreeSans 1200 0 0 0 io_in[29]
port 51 nsew
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 1200 0 0 0 io_in[2]
port 52 nsew
flabel metal3 s -960 371228 480 371468 0 FreeSans 1200 0 0 0 io_in[30]
port 53 nsew
flabel metal3 s -960 319140 480 319380 0 FreeSans 1200 0 0 0 io_in[31]
port 54 nsew
flabel metal3 s -960 267052 480 267292 0 FreeSans 1200 0 0 0 io_in[32]
port 55 nsew
flabel metal3 s -960 214828 480 215068 0 FreeSans 1200 0 0 0 io_in[33]
port 56 nsew
flabel metal3 s -960 162740 480 162980 0 FreeSans 1200 0 0 0 io_in[34]
port 57 nsew
flabel metal3 s -960 110516 480 110756 0 FreeSans 1200 0 0 0 io_in[35]
port 58 nsew
flabel metal3 s -960 71484 480 71724 0 FreeSans 1200 0 0 0 io_in[36]
port 59 nsew
flabel metal3 s -960 32316 480 32556 0 FreeSans 1200 0 0 0 io_in[37]
port 60 nsew
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 1200 0 0 0 io_in[3]
port 61 nsew
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 1200 0 0 0 io_in[4]
port 62 nsew
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 1200 0 0 0 io_in[5]
port 63 nsew
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 1200 0 0 0 io_in[6]
port 64 nsew
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 1200 0 0 0 io_in[7]
port 65 nsew
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 1200 0 0 0 io_in[8]
port 66 nsew
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 1200 0 0 0 io_in[9]
port 67 nsew
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 1200 0 0 0 io_oeb[0]
port 68 nsew
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 1200 0 0 0 io_oeb[10]
port 69 nsew
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 1200 0 0 0 io_oeb[11]
port 70 nsew
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 1200 0 0 0 io_oeb[12]
port 71 nsew
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 1200 0 0 0 io_oeb[13]
port 72 nsew
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 1200 0 0 0 io_oeb[14]
port 73 nsew
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 560 90 0 0 io_oeb[15]
port 74 nsew
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 560 90 0 0 io_oeb[16]
port 75 nsew
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 560 90 0 0 io_oeb[17]
port 76 nsew
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 560 90 0 0 io_oeb[18]
port 77 nsew
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 560 90 0 0 io_oeb[19]
port 78 nsew
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 1200 0 0 0 io_oeb[1]
port 79 nsew
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 560 90 0 0 io_oeb[20]
port 80 nsew
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 560 90 0 0 io_oeb[21]
port 81 nsew
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 560 90 0 0 io_oeb[22]
port 82 nsew
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 560 90 0 0 io_oeb[23]
port 83 nsew
flabel metal3 s -960 658052 480 658292 0 FreeSans 1200 0 0 0 io_oeb[24]
port 84 nsew
flabel metal3 s -960 605964 480 606204 0 FreeSans 1200 0 0 0 io_oeb[25]
port 85 nsew
flabel metal3 s -960 553740 480 553980 0 FreeSans 1200 0 0 0 io_oeb[26]
port 86 nsew
flabel metal3 s -960 501652 480 501892 0 FreeSans 1200 0 0 0 io_oeb[27]
port 87 nsew
flabel metal3 s -960 449428 480 449668 0 FreeSans 1200 0 0 0 io_oeb[28]
port 88 nsew
flabel metal3 s -960 397340 480 397580 0 FreeSans 1200 0 0 0 io_oeb[29]
port 89 nsew
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 1200 0 0 0 io_oeb[2]
port 90 nsew
flabel metal3 s -960 345252 480 345492 0 FreeSans 1200 0 0 0 io_oeb[30]
port 91 nsew
flabel metal3 s -960 293028 480 293268 0 FreeSans 1200 0 0 0 io_oeb[31]
port 92 nsew
flabel metal3 s -960 240940 480 241180 0 FreeSans 1200 0 0 0 io_oeb[32]
port 93 nsew
flabel metal3 s -960 188716 480 188956 0 FreeSans 1200 0 0 0 io_oeb[33]
port 94 nsew
flabel metal3 s -960 136628 480 136868 0 FreeSans 1200 0 0 0 io_oeb[34]
port 95 nsew
flabel metal3 s -960 84540 480 84780 0 FreeSans 1200 0 0 0 io_oeb[35]
port 96 nsew
flabel metal3 s -960 45372 480 45612 0 FreeSans 1200 0 0 0 io_oeb[36]
port 97 nsew
flabel metal3 s -960 6340 480 6580 0 FreeSans 1200 0 0 0 io_oeb[37]
port 98 nsew
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 1200 0 0 0 io_oeb[3]
port 99 nsew
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 1200 0 0 0 io_oeb[4]
port 100 nsew
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 1200 0 0 0 io_oeb[5]
port 101 nsew
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 1200 0 0 0 io_oeb[6]
port 102 nsew
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 1200 0 0 0 io_oeb[7]
port 103 nsew
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 1200 0 0 0 io_oeb[8]
port 104 nsew
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 1200 0 0 0 io_oeb[9]
port 105 nsew
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 1200 0 0 0 io_out[0]
port 106 nsew
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 1200 0 0 0 io_out[10]
port 107 nsew
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 1200 0 0 0 io_out[11]
port 108 nsew
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 1200 0 0 0 io_out[12]
port 109 nsew
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 1200 0 0 0 io_out[13]
port 110 nsew
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 1200 0 0 0 io_out[14]
port 111 nsew
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 560 90 0 0 io_out[15]
port 112 nsew
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 560 90 0 0 io_out[16]
port 113 nsew
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 560 90 0 0 io_out[17]
port 114 nsew
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 560 90 0 0 io_out[18]
port 115 nsew
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 560 90 0 0 io_out[19]
port 116 nsew
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 1200 0 0 0 io_out[1]
port 117 nsew
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 560 90 0 0 io_out[20]
port 118 nsew
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 560 90 0 0 io_out[21]
port 119 nsew
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 560 90 0 0 io_out[22]
port 120 nsew
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 560 90 0 0 io_out[23]
port 121 nsew
flabel metal3 s -960 671108 480 671348 0 FreeSans 1200 0 0 0 io_out[24]
port 122 nsew
flabel metal3 s -960 619020 480 619260 0 FreeSans 1200 0 0 0 io_out[25]
port 123 nsew
flabel metal3 s -960 566796 480 567036 0 FreeSans 1200 0 0 0 io_out[26]
port 124 nsew
flabel metal3 s -960 514708 480 514948 0 FreeSans 1200 0 0 0 io_out[27]
port 125 nsew
flabel metal3 s -960 462484 480 462724 0 FreeSans 1200 0 0 0 io_out[28]
port 126 nsew
flabel metal3 s -960 410396 480 410636 0 FreeSans 1200 0 0 0 io_out[29]
port 127 nsew
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 1200 0 0 0 io_out[2]
port 128 nsew
flabel metal3 s -960 358308 480 358548 0 FreeSans 1200 0 0 0 io_out[30]
port 129 nsew
flabel metal3 s -960 306084 480 306324 0 FreeSans 1200 0 0 0 io_out[31]
port 130 nsew
flabel metal3 s -960 253996 480 254236 0 FreeSans 1200 0 0 0 io_out[32]
port 131 nsew
flabel metal3 s -960 201772 480 202012 0 FreeSans 1200 0 0 0 io_out[33]
port 132 nsew
flabel metal3 s -960 149684 480 149924 0 FreeSans 1200 0 0 0 io_out[34]
port 133 nsew
flabel metal3 s -960 97460 480 97700 0 FreeSans 1200 0 0 0 io_out[35]
port 134 nsew
flabel metal3 s -960 58428 480 58668 0 FreeSans 1200 0 0 0 io_out[36]
port 135 nsew
flabel metal3 s -960 19260 480 19500 0 FreeSans 1200 0 0 0 io_out[37]
port 136 nsew
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 1200 0 0 0 io_out[3]
port 137 nsew
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 1200 0 0 0 io_out[4]
port 138 nsew
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 1200 0 0 0 io_out[5]
port 139 nsew
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 1200 0 0 0 io_out[6]
port 140 nsew
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 1200 0 0 0 io_out[7]
port 141 nsew
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 1200 0 0 0 io_out[8]
port 142 nsew
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 1200 0 0 0 io_out[9]
port 143 nsew
flabel metal2 s 125846 -960 125958 480 0 FreeSans 560 90 0 0 la_data_in[0]
port 144 nsew
flabel metal2 s 480506 -960 480618 480 0 FreeSans 560 90 0 0 la_data_in[100]
port 145 nsew
flabel metal2 s 484002 -960 484114 480 0 FreeSans 560 90 0 0 la_data_in[101]
port 146 nsew
flabel metal2 s 487590 -960 487702 480 0 FreeSans 560 90 0 0 la_data_in[102]
port 147 nsew
flabel metal2 s 491086 -960 491198 480 0 FreeSans 560 90 0 0 la_data_in[103]
port 148 nsew
flabel metal2 s 494674 -960 494786 480 0 FreeSans 560 90 0 0 la_data_in[104]
port 149 nsew
flabel metal2 s 498170 -960 498282 480 0 FreeSans 560 90 0 0 la_data_in[105]
port 150 nsew
flabel metal2 s 501758 -960 501870 480 0 FreeSans 560 90 0 0 la_data_in[106]
port 151 nsew
flabel metal2 s 505346 -960 505458 480 0 FreeSans 560 90 0 0 la_data_in[107]
port 152 nsew
flabel metal2 s 508842 -960 508954 480 0 FreeSans 560 90 0 0 la_data_in[108]
port 153 nsew
flabel metal2 s 512430 -960 512542 480 0 FreeSans 560 90 0 0 la_data_in[109]
port 154 nsew
flabel metal2 s 161266 -960 161378 480 0 FreeSans 560 90 0 0 la_data_in[10]
port 155 nsew
flabel metal2 s 515926 -960 516038 480 0 FreeSans 560 90 0 0 la_data_in[110]
port 156 nsew
flabel metal2 s 519514 -960 519626 480 0 FreeSans 560 90 0 0 la_data_in[111]
port 157 nsew
flabel metal2 s 523010 -960 523122 480 0 FreeSans 560 90 0 0 la_data_in[112]
port 158 nsew
flabel metal2 s 526598 -960 526710 480 0 FreeSans 560 90 0 0 la_data_in[113]
port 159 nsew
flabel metal2 s 530094 -960 530206 480 0 FreeSans 560 90 0 0 la_data_in[114]
port 160 nsew
flabel metal2 s 533682 -960 533794 480 0 FreeSans 560 90 0 0 la_data_in[115]
port 161 nsew
flabel metal2 s 537178 -960 537290 480 0 FreeSans 560 90 0 0 la_data_in[116]
port 162 nsew
flabel metal2 s 540766 -960 540878 480 0 FreeSans 560 90 0 0 la_data_in[117]
port 163 nsew
flabel metal2 s 544354 -960 544466 480 0 FreeSans 560 90 0 0 la_data_in[118]
port 164 nsew
flabel metal2 s 547850 -960 547962 480 0 FreeSans 560 90 0 0 la_data_in[119]
port 165 nsew
flabel metal2 s 164854 -960 164966 480 0 FreeSans 560 90 0 0 la_data_in[11]
port 166 nsew
flabel metal2 s 551438 -960 551550 480 0 FreeSans 560 90 0 0 la_data_in[120]
port 167 nsew
flabel metal2 s 554934 -960 555046 480 0 FreeSans 560 90 0 0 la_data_in[121]
port 168 nsew
flabel metal2 s 558522 -960 558634 480 0 FreeSans 560 90 0 0 la_data_in[122]
port 169 nsew
flabel metal2 s 562018 -960 562130 480 0 FreeSans 560 90 0 0 la_data_in[123]
port 170 nsew
flabel metal2 s 565606 -960 565718 480 0 FreeSans 560 90 0 0 la_data_in[124]
port 171 nsew
flabel metal2 s 569102 -960 569214 480 0 FreeSans 560 90 0 0 la_data_in[125]
port 172 nsew
flabel metal2 s 572690 -960 572802 480 0 FreeSans 560 90 0 0 la_data_in[126]
port 173 nsew
flabel metal2 s 576278 -960 576390 480 0 FreeSans 560 90 0 0 la_data_in[127]
port 174 nsew
flabel metal2 s 168350 -960 168462 480 0 FreeSans 560 90 0 0 la_data_in[12]
port 175 nsew
flabel metal2 s 171938 -960 172050 480 0 FreeSans 560 90 0 0 la_data_in[13]
port 176 nsew
flabel metal2 s 175434 -960 175546 480 0 FreeSans 560 90 0 0 la_data_in[14]
port 177 nsew
flabel metal2 s 179022 -960 179134 480 0 FreeSans 560 90 0 0 la_data_in[15]
port 178 nsew
flabel metal2 s 182518 -960 182630 480 0 FreeSans 560 90 0 0 la_data_in[16]
port 179 nsew
flabel metal2 s 186106 -960 186218 480 0 FreeSans 560 90 0 0 la_data_in[17]
port 180 nsew
flabel metal2 s 189694 -960 189806 480 0 FreeSans 560 90 0 0 la_data_in[18]
port 181 nsew
flabel metal2 s 193190 -960 193302 480 0 FreeSans 560 90 0 0 la_data_in[19]
port 182 nsew
flabel metal2 s 129342 -960 129454 480 0 FreeSans 560 90 0 0 la_data_in[1]
port 183 nsew
flabel metal2 s 196778 -960 196890 480 0 FreeSans 560 90 0 0 la_data_in[20]
port 184 nsew
flabel metal2 s 200274 -960 200386 480 0 FreeSans 560 90 0 0 la_data_in[21]
port 185 nsew
flabel metal2 s 203862 -960 203974 480 0 FreeSans 560 90 0 0 la_data_in[22]
port 186 nsew
flabel metal2 s 207358 -960 207470 480 0 FreeSans 560 90 0 0 la_data_in[23]
port 187 nsew
flabel metal2 s 210946 -960 211058 480 0 FreeSans 560 90 0 0 la_data_in[24]
port 188 nsew
flabel metal2 s 214442 -960 214554 480 0 FreeSans 560 90 0 0 la_data_in[25]
port 189 nsew
flabel metal2 s 218030 -960 218142 480 0 FreeSans 560 90 0 0 la_data_in[26]
port 190 nsew
flabel metal2 s 221526 -960 221638 480 0 FreeSans 560 90 0 0 la_data_in[27]
port 191 nsew
flabel metal2 s 225114 -960 225226 480 0 FreeSans 560 90 0 0 la_data_in[28]
port 192 nsew
flabel metal2 s 228702 -960 228814 480 0 FreeSans 560 90 0 0 la_data_in[29]
port 193 nsew
flabel metal2 s 132930 -960 133042 480 0 FreeSans 560 90 0 0 la_data_in[2]
port 194 nsew
flabel metal2 s 232198 -960 232310 480 0 FreeSans 560 90 0 0 la_data_in[30]
port 195 nsew
flabel metal2 s 235786 -960 235898 480 0 FreeSans 560 90 0 0 la_data_in[31]
port 196 nsew
flabel metal2 s 239282 -960 239394 480 0 FreeSans 560 90 0 0 la_data_in[32]
port 197 nsew
flabel metal2 s 242870 -960 242982 480 0 FreeSans 560 90 0 0 la_data_in[33]
port 198 nsew
flabel metal2 s 246366 -960 246478 480 0 FreeSans 560 90 0 0 la_data_in[34]
port 199 nsew
flabel metal2 s 249954 -960 250066 480 0 FreeSans 560 90 0 0 la_data_in[35]
port 200 nsew
flabel metal2 s 253450 -960 253562 480 0 FreeSans 560 90 0 0 la_data_in[36]
port 201 nsew
flabel metal2 s 257038 -960 257150 480 0 FreeSans 560 90 0 0 la_data_in[37]
port 202 nsew
flabel metal2 s 260626 -960 260738 480 0 FreeSans 560 90 0 0 la_data_in[38]
port 203 nsew
flabel metal2 s 264122 -960 264234 480 0 FreeSans 560 90 0 0 la_data_in[39]
port 204 nsew
flabel metal2 s 136426 -960 136538 480 0 FreeSans 560 90 0 0 la_data_in[3]
port 205 nsew
flabel metal2 s 267710 -960 267822 480 0 FreeSans 560 90 0 0 la_data_in[40]
port 206 nsew
flabel metal2 s 271206 -960 271318 480 0 FreeSans 560 90 0 0 la_data_in[41]
port 207 nsew
flabel metal2 s 274794 -960 274906 480 0 FreeSans 560 90 0 0 la_data_in[42]
port 208 nsew
flabel metal2 s 278290 -960 278402 480 0 FreeSans 560 90 0 0 la_data_in[43]
port 209 nsew
flabel metal2 s 281878 -960 281990 480 0 FreeSans 560 90 0 0 la_data_in[44]
port 210 nsew
flabel metal2 s 285374 -960 285486 480 0 FreeSans 560 90 0 0 la_data_in[45]
port 211 nsew
flabel metal2 s 288962 -960 289074 480 0 FreeSans 560 90 0 0 la_data_in[46]
port 212 nsew
flabel metal2 s 292550 -960 292662 480 0 FreeSans 560 90 0 0 la_data_in[47]
port 213 nsew
flabel metal2 s 296046 -960 296158 480 0 FreeSans 560 90 0 0 la_data_in[48]
port 214 nsew
flabel metal2 s 299634 -960 299746 480 0 FreeSans 560 90 0 0 la_data_in[49]
port 215 nsew
flabel metal2 s 140014 -960 140126 480 0 FreeSans 560 90 0 0 la_data_in[4]
port 216 nsew
flabel metal2 s 303130 -960 303242 480 0 FreeSans 560 90 0 0 la_data_in[50]
port 217 nsew
flabel metal2 s 306718 -960 306830 480 0 FreeSans 560 90 0 0 la_data_in[51]
port 218 nsew
flabel metal2 s 310214 -960 310326 480 0 FreeSans 560 90 0 0 la_data_in[52]
port 219 nsew
flabel metal2 s 313802 -960 313914 480 0 FreeSans 560 90 0 0 la_data_in[53]
port 220 nsew
flabel metal2 s 317298 -960 317410 480 0 FreeSans 560 90 0 0 la_data_in[54]
port 221 nsew
flabel metal2 s 320886 -960 320998 480 0 FreeSans 560 90 0 0 la_data_in[55]
port 222 nsew
flabel metal2 s 324382 -960 324494 480 0 FreeSans 560 90 0 0 la_data_in[56]
port 223 nsew
flabel metal2 s 327970 -960 328082 480 0 FreeSans 560 90 0 0 la_data_in[57]
port 224 nsew
flabel metal2 s 331558 -960 331670 480 0 FreeSans 560 90 0 0 la_data_in[58]
port 225 nsew
flabel metal2 s 335054 -960 335166 480 0 FreeSans 560 90 0 0 la_data_in[59]
port 226 nsew
flabel metal2 s 143510 -960 143622 480 0 FreeSans 560 90 0 0 la_data_in[5]
port 227 nsew
flabel metal2 s 338642 -960 338754 480 0 FreeSans 560 90 0 0 la_data_in[60]
port 228 nsew
flabel metal2 s 342138 -960 342250 480 0 FreeSans 560 90 0 0 la_data_in[61]
port 229 nsew
flabel metal2 s 345726 -960 345838 480 0 FreeSans 560 90 0 0 la_data_in[62]
port 230 nsew
flabel metal2 s 349222 -960 349334 480 0 FreeSans 560 90 0 0 la_data_in[63]
port 231 nsew
flabel metal2 s 352810 -960 352922 480 0 FreeSans 560 90 0 0 la_data_in[64]
port 232 nsew
flabel metal2 s 356306 -960 356418 480 0 FreeSans 560 90 0 0 la_data_in[65]
port 233 nsew
flabel metal2 s 359894 -960 360006 480 0 FreeSans 560 90 0 0 la_data_in[66]
port 234 nsew
flabel metal2 s 363482 -960 363594 480 0 FreeSans 560 90 0 0 la_data_in[67]
port 235 nsew
flabel metal2 s 366978 -960 367090 480 0 FreeSans 560 90 0 0 la_data_in[68]
port 236 nsew
flabel metal2 s 370566 -960 370678 480 0 FreeSans 560 90 0 0 la_data_in[69]
port 237 nsew
flabel metal2 s 147098 -960 147210 480 0 FreeSans 560 90 0 0 la_data_in[6]
port 238 nsew
flabel metal2 s 374062 -960 374174 480 0 FreeSans 560 90 0 0 la_data_in[70]
port 239 nsew
flabel metal2 s 377650 -960 377762 480 0 FreeSans 560 90 0 0 la_data_in[71]
port 240 nsew
flabel metal2 s 381146 -960 381258 480 0 FreeSans 560 90 0 0 la_data_in[72]
port 241 nsew
flabel metal2 s 384734 -960 384846 480 0 FreeSans 560 90 0 0 la_data_in[73]
port 242 nsew
flabel metal2 s 388230 -960 388342 480 0 FreeSans 560 90 0 0 la_data_in[74]
port 243 nsew
flabel metal2 s 391818 -960 391930 480 0 FreeSans 560 90 0 0 la_data_in[75]
port 244 nsew
flabel metal2 s 395314 -960 395426 480 0 FreeSans 560 90 0 0 la_data_in[76]
port 245 nsew
flabel metal2 s 398902 -960 399014 480 0 FreeSans 560 90 0 0 la_data_in[77]
port 246 nsew
flabel metal2 s 402490 -960 402602 480 0 FreeSans 560 90 0 0 la_data_in[78]
port 247 nsew
flabel metal2 s 405986 -960 406098 480 0 FreeSans 560 90 0 0 la_data_in[79]
port 248 nsew
flabel metal2 s 150594 -960 150706 480 0 FreeSans 560 90 0 0 la_data_in[7]
port 249 nsew
flabel metal2 s 409574 -960 409686 480 0 FreeSans 560 90 0 0 la_data_in[80]
port 250 nsew
flabel metal2 s 413070 -960 413182 480 0 FreeSans 560 90 0 0 la_data_in[81]
port 251 nsew
flabel metal2 s 416658 -960 416770 480 0 FreeSans 560 90 0 0 la_data_in[82]
port 252 nsew
flabel metal2 s 420154 -960 420266 480 0 FreeSans 560 90 0 0 la_data_in[83]
port 253 nsew
flabel metal2 s 423742 -960 423854 480 0 FreeSans 560 90 0 0 la_data_in[84]
port 254 nsew
flabel metal2 s 427238 -960 427350 480 0 FreeSans 560 90 0 0 la_data_in[85]
port 255 nsew
flabel metal2 s 430826 -960 430938 480 0 FreeSans 560 90 0 0 la_data_in[86]
port 256 nsew
flabel metal2 s 434414 -960 434526 480 0 FreeSans 560 90 0 0 la_data_in[87]
port 257 nsew
flabel metal2 s 437910 -960 438022 480 0 FreeSans 560 90 0 0 la_data_in[88]
port 258 nsew
flabel metal2 s 441498 -960 441610 480 0 FreeSans 560 90 0 0 la_data_in[89]
port 259 nsew
flabel metal2 s 154182 -960 154294 480 0 FreeSans 560 90 0 0 la_data_in[8]
port 260 nsew
flabel metal2 s 444994 -960 445106 480 0 FreeSans 560 90 0 0 la_data_in[90]
port 261 nsew
flabel metal2 s 448582 -960 448694 480 0 FreeSans 560 90 0 0 la_data_in[91]
port 262 nsew
flabel metal2 s 452078 -960 452190 480 0 FreeSans 560 90 0 0 la_data_in[92]
port 263 nsew
flabel metal2 s 455666 -960 455778 480 0 FreeSans 560 90 0 0 la_data_in[93]
port 264 nsew
flabel metal2 s 459162 -960 459274 480 0 FreeSans 560 90 0 0 la_data_in[94]
port 265 nsew
flabel metal2 s 462750 -960 462862 480 0 FreeSans 560 90 0 0 la_data_in[95]
port 266 nsew
flabel metal2 s 466246 -960 466358 480 0 FreeSans 560 90 0 0 la_data_in[96]
port 267 nsew
flabel metal2 s 469834 -960 469946 480 0 FreeSans 560 90 0 0 la_data_in[97]
port 268 nsew
flabel metal2 s 473422 -960 473534 480 0 FreeSans 560 90 0 0 la_data_in[98]
port 269 nsew
flabel metal2 s 476918 -960 477030 480 0 FreeSans 560 90 0 0 la_data_in[99]
port 270 nsew
flabel metal2 s 157770 -960 157882 480 0 FreeSans 560 90 0 0 la_data_in[9]
port 271 nsew
flabel metal2 s 126950 -960 127062 480 0 FreeSans 560 90 0 0 la_data_out[0]
port 272 nsew
flabel metal2 s 481702 -960 481814 480 0 FreeSans 560 90 0 0 la_data_out[100]
port 273 nsew
flabel metal2 s 485198 -960 485310 480 0 FreeSans 560 90 0 0 la_data_out[101]
port 274 nsew
flabel metal2 s 488786 -960 488898 480 0 FreeSans 560 90 0 0 la_data_out[102]
port 275 nsew
flabel metal2 s 492282 -960 492394 480 0 FreeSans 560 90 0 0 la_data_out[103]
port 276 nsew
flabel metal2 s 495870 -960 495982 480 0 FreeSans 560 90 0 0 la_data_out[104]
port 277 nsew
flabel metal2 s 499366 -960 499478 480 0 FreeSans 560 90 0 0 la_data_out[105]
port 278 nsew
flabel metal2 s 502954 -960 503066 480 0 FreeSans 560 90 0 0 la_data_out[106]
port 279 nsew
flabel metal2 s 506450 -960 506562 480 0 FreeSans 560 90 0 0 la_data_out[107]
port 280 nsew
flabel metal2 s 510038 -960 510150 480 0 FreeSans 560 90 0 0 la_data_out[108]
port 281 nsew
flabel metal2 s 513534 -960 513646 480 0 FreeSans 560 90 0 0 la_data_out[109]
port 282 nsew
flabel metal2 s 162462 -960 162574 480 0 FreeSans 560 90 0 0 la_data_out[10]
port 283 nsew
flabel metal2 s 517122 -960 517234 480 0 FreeSans 560 90 0 0 la_data_out[110]
port 284 nsew
flabel metal2 s 520710 -960 520822 480 0 FreeSans 560 90 0 0 la_data_out[111]
port 285 nsew
flabel metal2 s 524206 -960 524318 480 0 FreeSans 560 90 0 0 la_data_out[112]
port 286 nsew
flabel metal2 s 527794 -960 527906 480 0 FreeSans 560 90 0 0 la_data_out[113]
port 287 nsew
flabel metal2 s 531290 -960 531402 480 0 FreeSans 560 90 0 0 la_data_out[114]
port 288 nsew
flabel metal2 s 534878 -960 534990 480 0 FreeSans 560 90 0 0 la_data_out[115]
port 289 nsew
flabel metal2 s 538374 -960 538486 480 0 FreeSans 560 90 0 0 la_data_out[116]
port 290 nsew
flabel metal2 s 541962 -960 542074 480 0 FreeSans 560 90 0 0 la_data_out[117]
port 291 nsew
flabel metal2 s 545458 -960 545570 480 0 FreeSans 560 90 0 0 la_data_out[118]
port 292 nsew
flabel metal2 s 549046 -960 549158 480 0 FreeSans 560 90 0 0 la_data_out[119]
port 293 nsew
flabel metal2 s 166050 -960 166162 480 0 FreeSans 560 90 0 0 la_data_out[11]
port 294 nsew
flabel metal2 s 552634 -960 552746 480 0 FreeSans 560 90 0 0 la_data_out[120]
port 295 nsew
flabel metal2 s 556130 -960 556242 480 0 FreeSans 560 90 0 0 la_data_out[121]
port 296 nsew
flabel metal2 s 559718 -960 559830 480 0 FreeSans 560 90 0 0 la_data_out[122]
port 297 nsew
flabel metal2 s 563214 -960 563326 480 0 FreeSans 560 90 0 0 la_data_out[123]
port 298 nsew
flabel metal2 s 566802 -960 566914 480 0 FreeSans 560 90 0 0 la_data_out[124]
port 299 nsew
flabel metal2 s 570298 -960 570410 480 0 FreeSans 560 90 0 0 la_data_out[125]
port 300 nsew
flabel metal2 s 573886 -960 573998 480 0 FreeSans 560 90 0 0 la_data_out[126]
port 301 nsew
flabel metal2 s 577382 -960 577494 480 0 FreeSans 560 90 0 0 la_data_out[127]
port 302 nsew
flabel metal2 s 169546 -960 169658 480 0 FreeSans 560 90 0 0 la_data_out[12]
port 303 nsew
flabel metal2 s 173134 -960 173246 480 0 FreeSans 560 90 0 0 la_data_out[13]
port 304 nsew
flabel metal2 s 176630 -960 176742 480 0 FreeSans 560 90 0 0 la_data_out[14]
port 305 nsew
flabel metal2 s 180218 -960 180330 480 0 FreeSans 560 90 0 0 la_data_out[15]
port 306 nsew
flabel metal2 s 183714 -960 183826 480 0 FreeSans 560 90 0 0 la_data_out[16]
port 307 nsew
flabel metal2 s 187302 -960 187414 480 0 FreeSans 560 90 0 0 la_data_out[17]
port 308 nsew
flabel metal2 s 190798 -960 190910 480 0 FreeSans 560 90 0 0 la_data_out[18]
port 309 nsew
flabel metal2 s 194386 -960 194498 480 0 FreeSans 560 90 0 0 la_data_out[19]
port 310 nsew
flabel metal2 s 130538 -960 130650 480 0 FreeSans 560 90 0 0 la_data_out[1]
port 311 nsew
flabel metal2 s 197882 -960 197994 480 0 FreeSans 560 90 0 0 la_data_out[20]
port 312 nsew
flabel metal2 s 201470 -960 201582 480 0 FreeSans 560 90 0 0 la_data_out[21]
port 313 nsew
flabel metal2 s 205058 -960 205170 480 0 FreeSans 560 90 0 0 la_data_out[22]
port 314 nsew
flabel metal2 s 208554 -960 208666 480 0 FreeSans 560 90 0 0 la_data_out[23]
port 315 nsew
flabel metal2 s 212142 -960 212254 480 0 FreeSans 560 90 0 0 la_data_out[24]
port 316 nsew
flabel metal2 s 215638 -960 215750 480 0 FreeSans 560 90 0 0 la_data_out[25]
port 317 nsew
flabel metal2 s 219226 -960 219338 480 0 FreeSans 560 90 0 0 la_data_out[26]
port 318 nsew
flabel metal2 s 222722 -960 222834 480 0 FreeSans 560 90 0 0 la_data_out[27]
port 319 nsew
flabel metal2 s 226310 -960 226422 480 0 FreeSans 560 90 0 0 la_data_out[28]
port 320 nsew
flabel metal2 s 229806 -960 229918 480 0 FreeSans 560 90 0 0 la_data_out[29]
port 321 nsew
flabel metal2 s 134126 -960 134238 480 0 FreeSans 560 90 0 0 la_data_out[2]
port 322 nsew
flabel metal2 s 233394 -960 233506 480 0 FreeSans 560 90 0 0 la_data_out[30]
port 323 nsew
flabel metal2 s 236982 -960 237094 480 0 FreeSans 560 90 0 0 la_data_out[31]
port 324 nsew
flabel metal2 s 240478 -960 240590 480 0 FreeSans 560 90 0 0 la_data_out[32]
port 325 nsew
flabel metal2 s 244066 -960 244178 480 0 FreeSans 560 90 0 0 la_data_out[33]
port 326 nsew
flabel metal2 s 247562 -960 247674 480 0 FreeSans 560 90 0 0 la_data_out[34]
port 327 nsew
flabel metal2 s 251150 -960 251262 480 0 FreeSans 560 90 0 0 la_data_out[35]
port 328 nsew
flabel metal2 s 254646 -960 254758 480 0 FreeSans 560 90 0 0 la_data_out[36]
port 329 nsew
flabel metal2 s 258234 -960 258346 480 0 FreeSans 560 90 0 0 la_data_out[37]
port 330 nsew
flabel metal2 s 261730 -960 261842 480 0 FreeSans 560 90 0 0 la_data_out[38]
port 331 nsew
flabel metal2 s 265318 -960 265430 480 0 FreeSans 560 90 0 0 la_data_out[39]
port 332 nsew
flabel metal2 s 137622 -960 137734 480 0 FreeSans 560 90 0 0 la_data_out[3]
port 333 nsew
flabel metal2 s 268814 -960 268926 480 0 FreeSans 560 90 0 0 la_data_out[40]
port 334 nsew
flabel metal2 s 272402 -960 272514 480 0 FreeSans 560 90 0 0 la_data_out[41]
port 335 nsew
flabel metal2 s 275990 -960 276102 480 0 FreeSans 560 90 0 0 la_data_out[42]
port 336 nsew
flabel metal2 s 279486 -960 279598 480 0 FreeSans 560 90 0 0 la_data_out[43]
port 337 nsew
flabel metal2 s 283074 -960 283186 480 0 FreeSans 560 90 0 0 la_data_out[44]
port 338 nsew
flabel metal2 s 286570 -960 286682 480 0 FreeSans 560 90 0 0 la_data_out[45]
port 339 nsew
flabel metal2 s 290158 -960 290270 480 0 FreeSans 560 90 0 0 la_data_out[46]
port 340 nsew
flabel metal2 s 293654 -960 293766 480 0 FreeSans 560 90 0 0 la_data_out[47]
port 341 nsew
flabel metal2 s 297242 -960 297354 480 0 FreeSans 560 90 0 0 la_data_out[48]
port 342 nsew
flabel metal2 s 300738 -960 300850 480 0 FreeSans 560 90 0 0 la_data_out[49]
port 343 nsew
flabel metal2 s 141210 -960 141322 480 0 FreeSans 560 90 0 0 la_data_out[4]
port 344 nsew
flabel metal2 s 304326 -960 304438 480 0 FreeSans 560 90 0 0 la_data_out[50]
port 345 nsew
flabel metal2 s 307914 -960 308026 480 0 FreeSans 560 90 0 0 la_data_out[51]
port 346 nsew
flabel metal2 s 311410 -960 311522 480 0 FreeSans 560 90 0 0 la_data_out[52]
port 347 nsew
flabel metal2 s 314998 -960 315110 480 0 FreeSans 560 90 0 0 la_data_out[53]
port 348 nsew
flabel metal2 s 318494 -960 318606 480 0 FreeSans 560 90 0 0 la_data_out[54]
port 349 nsew
flabel metal2 s 322082 -960 322194 480 0 FreeSans 560 90 0 0 la_data_out[55]
port 350 nsew
flabel metal2 s 325578 -960 325690 480 0 FreeSans 560 90 0 0 la_data_out[56]
port 351 nsew
flabel metal2 s 329166 -960 329278 480 0 FreeSans 560 90 0 0 la_data_out[57]
port 352 nsew
flabel metal2 s 332662 -960 332774 480 0 FreeSans 560 90 0 0 la_data_out[58]
port 353 nsew
flabel metal2 s 336250 -960 336362 480 0 FreeSans 560 90 0 0 la_data_out[59]
port 354 nsew
flabel metal2 s 144706 -960 144818 480 0 FreeSans 560 90 0 0 la_data_out[5]
port 355 nsew
flabel metal2 s 339838 -960 339950 480 0 FreeSans 560 90 0 0 la_data_out[60]
port 356 nsew
flabel metal2 s 343334 -960 343446 480 0 FreeSans 560 90 0 0 la_data_out[61]
port 357 nsew
flabel metal2 s 346922 -960 347034 480 0 FreeSans 560 90 0 0 la_data_out[62]
port 358 nsew
flabel metal2 s 350418 -960 350530 480 0 FreeSans 560 90 0 0 la_data_out[63]
port 359 nsew
flabel metal2 s 354006 -960 354118 480 0 FreeSans 560 90 0 0 la_data_out[64]
port 360 nsew
flabel metal2 s 357502 -960 357614 480 0 FreeSans 560 90 0 0 la_data_out[65]
port 361 nsew
flabel metal2 s 361090 -960 361202 480 0 FreeSans 560 90 0 0 la_data_out[66]
port 362 nsew
flabel metal2 s 364586 -960 364698 480 0 FreeSans 560 90 0 0 la_data_out[67]
port 363 nsew
flabel metal2 s 368174 -960 368286 480 0 FreeSans 560 90 0 0 la_data_out[68]
port 364 nsew
flabel metal2 s 371670 -960 371782 480 0 FreeSans 560 90 0 0 la_data_out[69]
port 365 nsew
flabel metal2 s 148294 -960 148406 480 0 FreeSans 560 90 0 0 la_data_out[6]
port 366 nsew
flabel metal2 s 375258 -960 375370 480 0 FreeSans 560 90 0 0 la_data_out[70]
port 367 nsew
flabel metal2 s 378846 -960 378958 480 0 FreeSans 560 90 0 0 la_data_out[71]
port 368 nsew
flabel metal2 s 382342 -960 382454 480 0 FreeSans 560 90 0 0 la_data_out[72]
port 369 nsew
flabel metal2 s 385930 -960 386042 480 0 FreeSans 560 90 0 0 la_data_out[73]
port 370 nsew
flabel metal2 s 389426 -960 389538 480 0 FreeSans 560 90 0 0 la_data_out[74]
port 371 nsew
flabel metal2 s 393014 -960 393126 480 0 FreeSans 560 90 0 0 la_data_out[75]
port 372 nsew
flabel metal2 s 396510 -960 396622 480 0 FreeSans 560 90 0 0 la_data_out[76]
port 373 nsew
flabel metal2 s 400098 -960 400210 480 0 FreeSans 560 90 0 0 la_data_out[77]
port 374 nsew
flabel metal2 s 403594 -960 403706 480 0 FreeSans 560 90 0 0 la_data_out[78]
port 375 nsew
flabel metal2 s 407182 -960 407294 480 0 FreeSans 560 90 0 0 la_data_out[79]
port 376 nsew
flabel metal2 s 151790 -960 151902 480 0 FreeSans 560 90 0 0 la_data_out[7]
port 377 nsew
flabel metal2 s 410770 -960 410882 480 0 FreeSans 560 90 0 0 la_data_out[80]
port 378 nsew
flabel metal2 s 414266 -960 414378 480 0 FreeSans 560 90 0 0 la_data_out[81]
port 379 nsew
flabel metal2 s 417854 -960 417966 480 0 FreeSans 560 90 0 0 la_data_out[82]
port 380 nsew
flabel metal2 s 421350 -960 421462 480 0 FreeSans 560 90 0 0 la_data_out[83]
port 381 nsew
flabel metal2 s 424938 -960 425050 480 0 FreeSans 560 90 0 0 la_data_out[84]
port 382 nsew
flabel metal2 s 428434 -960 428546 480 0 FreeSans 560 90 0 0 la_data_out[85]
port 383 nsew
flabel metal2 s 432022 -960 432134 480 0 FreeSans 560 90 0 0 la_data_out[86]
port 384 nsew
flabel metal2 s 435518 -960 435630 480 0 FreeSans 560 90 0 0 la_data_out[87]
port 385 nsew
flabel metal2 s 439106 -960 439218 480 0 FreeSans 560 90 0 0 la_data_out[88]
port 386 nsew
flabel metal2 s 442602 -960 442714 480 0 FreeSans 560 90 0 0 la_data_out[89]
port 387 nsew
flabel metal2 s 155378 -960 155490 480 0 FreeSans 560 90 0 0 la_data_out[8]
port 388 nsew
flabel metal2 s 446190 -960 446302 480 0 FreeSans 560 90 0 0 la_data_out[90]
port 389 nsew
flabel metal2 s 449778 -960 449890 480 0 FreeSans 560 90 0 0 la_data_out[91]
port 390 nsew
flabel metal2 s 453274 -960 453386 480 0 FreeSans 560 90 0 0 la_data_out[92]
port 391 nsew
flabel metal2 s 456862 -960 456974 480 0 FreeSans 560 90 0 0 la_data_out[93]
port 392 nsew
flabel metal2 s 460358 -960 460470 480 0 FreeSans 560 90 0 0 la_data_out[94]
port 393 nsew
flabel metal2 s 463946 -960 464058 480 0 FreeSans 560 90 0 0 la_data_out[95]
port 394 nsew
flabel metal2 s 467442 -960 467554 480 0 FreeSans 560 90 0 0 la_data_out[96]
port 395 nsew
flabel metal2 s 471030 -960 471142 480 0 FreeSans 560 90 0 0 la_data_out[97]
port 396 nsew
flabel metal2 s 474526 -960 474638 480 0 FreeSans 560 90 0 0 la_data_out[98]
port 397 nsew
flabel metal2 s 478114 -960 478226 480 0 FreeSans 560 90 0 0 la_data_out[99]
port 398 nsew
flabel metal2 s 158874 -960 158986 480 0 FreeSans 560 90 0 0 la_data_out[9]
port 399 nsew
flabel metal2 s 128146 -960 128258 480 0 FreeSans 560 90 0 0 la_oenb[0]
port 400 nsew
flabel metal2 s 482806 -960 482918 480 0 FreeSans 560 90 0 0 la_oenb[100]
port 401 nsew
flabel metal2 s 486394 -960 486506 480 0 FreeSans 560 90 0 0 la_oenb[101]
port 402 nsew
flabel metal2 s 489890 -960 490002 480 0 FreeSans 560 90 0 0 la_oenb[102]
port 403 nsew
flabel metal2 s 493478 -960 493590 480 0 FreeSans 560 90 0 0 la_oenb[103]
port 404 nsew
flabel metal2 s 497066 -960 497178 480 0 FreeSans 560 90 0 0 la_oenb[104]
port 405 nsew
flabel metal2 s 500562 -960 500674 480 0 FreeSans 560 90 0 0 la_oenb[105]
port 406 nsew
flabel metal2 s 504150 -960 504262 480 0 FreeSans 560 90 0 0 la_oenb[106]
port 407 nsew
flabel metal2 s 507646 -960 507758 480 0 FreeSans 560 90 0 0 la_oenb[107]
port 408 nsew
flabel metal2 s 511234 -960 511346 480 0 FreeSans 560 90 0 0 la_oenb[108]
port 409 nsew
flabel metal2 s 514730 -960 514842 480 0 FreeSans 560 90 0 0 la_oenb[109]
port 410 nsew
flabel metal2 s 163658 -960 163770 480 0 FreeSans 560 90 0 0 la_oenb[10]
port 411 nsew
flabel metal2 s 518318 -960 518430 480 0 FreeSans 560 90 0 0 la_oenb[110]
port 412 nsew
flabel metal2 s 521814 -960 521926 480 0 FreeSans 560 90 0 0 la_oenb[111]
port 413 nsew
flabel metal2 s 525402 -960 525514 480 0 FreeSans 560 90 0 0 la_oenb[112]
port 414 nsew
flabel metal2 s 528990 -960 529102 480 0 FreeSans 560 90 0 0 la_oenb[113]
port 415 nsew
flabel metal2 s 532486 -960 532598 480 0 FreeSans 560 90 0 0 la_oenb[114]
port 416 nsew
flabel metal2 s 536074 -960 536186 480 0 FreeSans 560 90 0 0 la_oenb[115]
port 417 nsew
flabel metal2 s 539570 -960 539682 480 0 FreeSans 560 90 0 0 la_oenb[116]
port 418 nsew
flabel metal2 s 543158 -960 543270 480 0 FreeSans 560 90 0 0 la_oenb[117]
port 419 nsew
flabel metal2 s 546654 -960 546766 480 0 FreeSans 560 90 0 0 la_oenb[118]
port 420 nsew
flabel metal2 s 550242 -960 550354 480 0 FreeSans 560 90 0 0 la_oenb[119]
port 421 nsew
flabel metal2 s 167154 -960 167266 480 0 FreeSans 560 90 0 0 la_oenb[11]
port 422 nsew
flabel metal2 s 553738 -960 553850 480 0 FreeSans 560 90 0 0 la_oenb[120]
port 423 nsew
flabel metal2 s 557326 -960 557438 480 0 FreeSans 560 90 0 0 la_oenb[121]
port 424 nsew
flabel metal2 s 560822 -960 560934 480 0 FreeSans 560 90 0 0 la_oenb[122]
port 425 nsew
flabel metal2 s 564410 -960 564522 480 0 FreeSans 560 90 0 0 la_oenb[123]
port 426 nsew
flabel metal2 s 567998 -960 568110 480 0 FreeSans 560 90 0 0 la_oenb[124]
port 427 nsew
flabel metal2 s 571494 -960 571606 480 0 FreeSans 560 90 0 0 la_oenb[125]
port 428 nsew
flabel metal2 s 575082 -960 575194 480 0 FreeSans 560 90 0 0 la_oenb[126]
port 429 nsew
flabel metal2 s 578578 -960 578690 480 0 FreeSans 560 90 0 0 la_oenb[127]
port 430 nsew
flabel metal2 s 170742 -960 170854 480 0 FreeSans 560 90 0 0 la_oenb[12]
port 431 nsew
flabel metal2 s 174238 -960 174350 480 0 FreeSans 560 90 0 0 la_oenb[13]
port 432 nsew
flabel metal2 s 177826 -960 177938 480 0 FreeSans 560 90 0 0 la_oenb[14]
port 433 nsew
flabel metal2 s 181414 -960 181526 480 0 FreeSans 560 90 0 0 la_oenb[15]
port 434 nsew
flabel metal2 s 184910 -960 185022 480 0 FreeSans 560 90 0 0 la_oenb[16]
port 435 nsew
flabel metal2 s 188498 -960 188610 480 0 FreeSans 560 90 0 0 la_oenb[17]
port 436 nsew
flabel metal2 s 191994 -960 192106 480 0 FreeSans 560 90 0 0 la_oenb[18]
port 437 nsew
flabel metal2 s 195582 -960 195694 480 0 FreeSans 560 90 0 0 la_oenb[19]
port 438 nsew
flabel metal2 s 131734 -960 131846 480 0 FreeSans 560 90 0 0 la_oenb[1]
port 439 nsew
flabel metal2 s 199078 -960 199190 480 0 FreeSans 560 90 0 0 la_oenb[20]
port 440 nsew
flabel metal2 s 202666 -960 202778 480 0 FreeSans 560 90 0 0 la_oenb[21]
port 441 nsew
flabel metal2 s 206162 -960 206274 480 0 FreeSans 560 90 0 0 la_oenb[22]
port 442 nsew
flabel metal2 s 209750 -960 209862 480 0 FreeSans 560 90 0 0 la_oenb[23]
port 443 nsew
flabel metal2 s 213338 -960 213450 480 0 FreeSans 560 90 0 0 la_oenb[24]
port 444 nsew
flabel metal2 s 216834 -960 216946 480 0 FreeSans 560 90 0 0 la_oenb[25]
port 445 nsew
flabel metal2 s 220422 -960 220534 480 0 FreeSans 560 90 0 0 la_oenb[26]
port 446 nsew
flabel metal2 s 223918 -960 224030 480 0 FreeSans 560 90 0 0 la_oenb[27]
port 447 nsew
flabel metal2 s 227506 -960 227618 480 0 FreeSans 560 90 0 0 la_oenb[28]
port 448 nsew
flabel metal2 s 231002 -960 231114 480 0 FreeSans 560 90 0 0 la_oenb[29]
port 449 nsew
flabel metal2 s 135230 -960 135342 480 0 FreeSans 560 90 0 0 la_oenb[2]
port 450 nsew
flabel metal2 s 234590 -960 234702 480 0 FreeSans 560 90 0 0 la_oenb[30]
port 451 nsew
flabel metal2 s 238086 -960 238198 480 0 FreeSans 560 90 0 0 la_oenb[31]
port 452 nsew
flabel metal2 s 241674 -960 241786 480 0 FreeSans 560 90 0 0 la_oenb[32]
port 453 nsew
flabel metal2 s 245170 -960 245282 480 0 FreeSans 560 90 0 0 la_oenb[33]
port 454 nsew
flabel metal2 s 248758 -960 248870 480 0 FreeSans 560 90 0 0 la_oenb[34]
port 455 nsew
flabel metal2 s 252346 -960 252458 480 0 FreeSans 560 90 0 0 la_oenb[35]
port 456 nsew
flabel metal2 s 255842 -960 255954 480 0 FreeSans 560 90 0 0 la_oenb[36]
port 457 nsew
flabel metal2 s 259430 -960 259542 480 0 FreeSans 560 90 0 0 la_oenb[37]
port 458 nsew
flabel metal2 s 262926 -960 263038 480 0 FreeSans 560 90 0 0 la_oenb[38]
port 459 nsew
flabel metal2 s 266514 -960 266626 480 0 FreeSans 560 90 0 0 la_oenb[39]
port 460 nsew
flabel metal2 s 138818 -960 138930 480 0 FreeSans 560 90 0 0 la_oenb[3]
port 461 nsew
flabel metal2 s 270010 -960 270122 480 0 FreeSans 560 90 0 0 la_oenb[40]
port 462 nsew
flabel metal2 s 273598 -960 273710 480 0 FreeSans 560 90 0 0 la_oenb[41]
port 463 nsew
flabel metal2 s 277094 -960 277206 480 0 FreeSans 560 90 0 0 la_oenb[42]
port 464 nsew
flabel metal2 s 280682 -960 280794 480 0 FreeSans 560 90 0 0 la_oenb[43]
port 465 nsew
flabel metal2 s 284270 -960 284382 480 0 FreeSans 560 90 0 0 la_oenb[44]
port 466 nsew
flabel metal2 s 287766 -960 287878 480 0 FreeSans 560 90 0 0 la_oenb[45]
port 467 nsew
flabel metal2 s 291354 -960 291466 480 0 FreeSans 560 90 0 0 la_oenb[46]
port 468 nsew
flabel metal2 s 294850 -960 294962 480 0 FreeSans 560 90 0 0 la_oenb[47]
port 469 nsew
flabel metal2 s 298438 -960 298550 480 0 FreeSans 560 90 0 0 la_oenb[48]
port 470 nsew
flabel metal2 s 301934 -960 302046 480 0 FreeSans 560 90 0 0 la_oenb[49]
port 471 nsew
flabel metal2 s 142406 -960 142518 480 0 FreeSans 560 90 0 0 la_oenb[4]
port 472 nsew
flabel metal2 s 305522 -960 305634 480 0 FreeSans 560 90 0 0 la_oenb[50]
port 473 nsew
flabel metal2 s 309018 -960 309130 480 0 FreeSans 560 90 0 0 la_oenb[51]
port 474 nsew
flabel metal2 s 312606 -960 312718 480 0 FreeSans 560 90 0 0 la_oenb[52]
port 475 nsew
flabel metal2 s 316194 -960 316306 480 0 FreeSans 560 90 0 0 la_oenb[53]
port 476 nsew
flabel metal2 s 319690 -960 319802 480 0 FreeSans 560 90 0 0 la_oenb[54]
port 477 nsew
flabel metal2 s 323278 -960 323390 480 0 FreeSans 560 90 0 0 la_oenb[55]
port 478 nsew
flabel metal2 s 326774 -960 326886 480 0 FreeSans 560 90 0 0 la_oenb[56]
port 479 nsew
flabel metal2 s 330362 -960 330474 480 0 FreeSans 560 90 0 0 la_oenb[57]
port 480 nsew
flabel metal2 s 333858 -960 333970 480 0 FreeSans 560 90 0 0 la_oenb[58]
port 481 nsew
flabel metal2 s 337446 -960 337558 480 0 FreeSans 560 90 0 0 la_oenb[59]
port 482 nsew
flabel metal2 s 145902 -960 146014 480 0 FreeSans 560 90 0 0 la_oenb[5]
port 483 nsew
flabel metal2 s 340942 -960 341054 480 0 FreeSans 560 90 0 0 la_oenb[60]
port 484 nsew
flabel metal2 s 344530 -960 344642 480 0 FreeSans 560 90 0 0 la_oenb[61]
port 485 nsew
flabel metal2 s 348026 -960 348138 480 0 FreeSans 560 90 0 0 la_oenb[62]
port 486 nsew
flabel metal2 s 351614 -960 351726 480 0 FreeSans 560 90 0 0 la_oenb[63]
port 487 nsew
flabel metal2 s 355202 -960 355314 480 0 FreeSans 560 90 0 0 la_oenb[64]
port 488 nsew
flabel metal2 s 358698 -960 358810 480 0 FreeSans 560 90 0 0 la_oenb[65]
port 489 nsew
flabel metal2 s 362286 -960 362398 480 0 FreeSans 560 90 0 0 la_oenb[66]
port 490 nsew
flabel metal2 s 365782 -960 365894 480 0 FreeSans 560 90 0 0 la_oenb[67]
port 491 nsew
flabel metal2 s 369370 -960 369482 480 0 FreeSans 560 90 0 0 la_oenb[68]
port 492 nsew
flabel metal2 s 372866 -960 372978 480 0 FreeSans 560 90 0 0 la_oenb[69]
port 493 nsew
flabel metal2 s 149490 -960 149602 480 0 FreeSans 560 90 0 0 la_oenb[6]
port 494 nsew
flabel metal2 s 376454 -960 376566 480 0 FreeSans 560 90 0 0 la_oenb[70]
port 495 nsew
flabel metal2 s 379950 -960 380062 480 0 FreeSans 560 90 0 0 la_oenb[71]
port 496 nsew
flabel metal2 s 383538 -960 383650 480 0 FreeSans 560 90 0 0 la_oenb[72]
port 497 nsew
flabel metal2 s 387126 -960 387238 480 0 FreeSans 560 90 0 0 la_oenb[73]
port 498 nsew
flabel metal2 s 390622 -960 390734 480 0 FreeSans 560 90 0 0 la_oenb[74]
port 499 nsew
flabel metal2 s 394210 -960 394322 480 0 FreeSans 560 90 0 0 la_oenb[75]
port 500 nsew
flabel metal2 s 397706 -960 397818 480 0 FreeSans 560 90 0 0 la_oenb[76]
port 501 nsew
flabel metal2 s 401294 -960 401406 480 0 FreeSans 560 90 0 0 la_oenb[77]
port 502 nsew
flabel metal2 s 404790 -960 404902 480 0 FreeSans 560 90 0 0 la_oenb[78]
port 503 nsew
flabel metal2 s 408378 -960 408490 480 0 FreeSans 560 90 0 0 la_oenb[79]
port 504 nsew
flabel metal2 s 152986 -960 153098 480 0 FreeSans 560 90 0 0 la_oenb[7]
port 505 nsew
flabel metal2 s 411874 -960 411986 480 0 FreeSans 560 90 0 0 la_oenb[80]
port 506 nsew
flabel metal2 s 415462 -960 415574 480 0 FreeSans 560 90 0 0 la_oenb[81]
port 507 nsew
flabel metal2 s 418958 -960 419070 480 0 FreeSans 560 90 0 0 la_oenb[82]
port 508 nsew
flabel metal2 s 422546 -960 422658 480 0 FreeSans 560 90 0 0 la_oenb[83]
port 509 nsew
flabel metal2 s 426134 -960 426246 480 0 FreeSans 560 90 0 0 la_oenb[84]
port 510 nsew
flabel metal2 s 429630 -960 429742 480 0 FreeSans 560 90 0 0 la_oenb[85]
port 511 nsew
flabel metal2 s 433218 -960 433330 480 0 FreeSans 560 90 0 0 la_oenb[86]
port 512 nsew
flabel metal2 s 436714 -960 436826 480 0 FreeSans 560 90 0 0 la_oenb[87]
port 513 nsew
flabel metal2 s 440302 -960 440414 480 0 FreeSans 560 90 0 0 la_oenb[88]
port 514 nsew
flabel metal2 s 443798 -960 443910 480 0 FreeSans 560 90 0 0 la_oenb[89]
port 515 nsew
flabel metal2 s 156574 -960 156686 480 0 FreeSans 560 90 0 0 la_oenb[8]
port 516 nsew
flabel metal2 s 447386 -960 447498 480 0 FreeSans 560 90 0 0 la_oenb[90]
port 517 nsew
flabel metal2 s 450882 -960 450994 480 0 FreeSans 560 90 0 0 la_oenb[91]
port 518 nsew
flabel metal2 s 454470 -960 454582 480 0 FreeSans 560 90 0 0 la_oenb[92]
port 519 nsew
flabel metal2 s 458058 -960 458170 480 0 FreeSans 560 90 0 0 la_oenb[93]
port 520 nsew
flabel metal2 s 461554 -960 461666 480 0 FreeSans 560 90 0 0 la_oenb[94]
port 521 nsew
flabel metal2 s 465142 -960 465254 480 0 FreeSans 560 90 0 0 la_oenb[95]
port 522 nsew
flabel metal2 s 468638 -960 468750 480 0 FreeSans 560 90 0 0 la_oenb[96]
port 523 nsew
flabel metal2 s 472226 -960 472338 480 0 FreeSans 560 90 0 0 la_oenb[97]
port 524 nsew
flabel metal2 s 475722 -960 475834 480 0 FreeSans 560 90 0 0 la_oenb[98]
port 525 nsew
flabel metal2 s 479310 -960 479422 480 0 FreeSans 560 90 0 0 la_oenb[99]
port 526 nsew
flabel metal2 s 160070 -960 160182 480 0 FreeSans 560 90 0 0 la_oenb[9]
port 527 nsew
flabel metal2 s 579774 -960 579886 480 0 FreeSans 560 90 0 0 user_clock2
port 528 nsew
flabel metal2 s 580970 -960 581082 480 0 FreeSans 560 90 0 0 user_irq[0]
port 529 nsew
flabel metal2 s 582166 -960 582278 480 0 FreeSans 560 90 0 0 user_irq[1]
port 530 nsew
flabel metal2 s 583362 -960 583474 480 0 FreeSans 560 90 0 0 user_irq[2]
port 531 nsew
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 73794 -7654 74414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 109794 -7654 110414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 145794 -7654 146414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 181794 -7654 182414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 217794 -7654 218414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 253794 -7654 254414 4103 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 253794 27193 254414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 289794 -7654 290414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 45234 -7654 45854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 81234 -7654 81854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 117234 -7654 117854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 153234 -7654 153854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 189234 -7654 189854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 225234 -7654 225854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 261234 -7654 261854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 297234 -7654 297854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 333234 -7654 333854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 369234 354900 369854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 405234 -7654 405854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 441234 -7654 441854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 477234 354900 477854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 513234 -7654 513854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 549234 -7654 549854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 16674 -7654 17294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 52674 -7654 53294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 88674 -7654 89294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 124674 -7654 125294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 160674 -7654 161294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 196674 -7654 197294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 232674 -7654 233294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 268674 -7654 269294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 304674 -7654 305294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 340674 -7654 341294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 376674 -7654 377294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 412674 -7654 413294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 448674 -7654 449294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 484674 -7654 485294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 520674 -7654 521294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 556674 -7654 557294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 24114 -7654 24734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 60114 -7654 60734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 96114 -7654 96734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 132114 -7654 132734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 168114 -7654 168734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 204114 -7654 204734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 240114 27193 240734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 276114 -7654 276734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 312114 -7654 312734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 348114 -7654 348734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 384114 -7654 384734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 420114 -7654 420734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 456114 -7654 456734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 492114 354900 492734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 528114 -7654 528734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 564114 -7654 564734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 20394 -7654 21014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 56394 -7654 57014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 92394 354900 93014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 128394 -7654 129014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 164394 -7654 165014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 200394 354900 201014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 236394 -7654 237014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 272394 -7654 273014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 308394 354900 309014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 344394 -7654 345014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 380394 -7654 381014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 416394 -7654 417014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 452394 -7654 453014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 488394 -7654 489014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 524394 -7654 525014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 560394 -7654 561014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 27834 -7654 28454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 63834 -7654 64454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 99834 -7654 100454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 135834 -7654 136454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 171834 -7654 172454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 207834 -7654 208454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 243834 27193 244454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 279834 -7654 280454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 315834 -7654 316454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 351834 -7654 352454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 387834 -7654 388454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 423834 -7654 424454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 459834 -7654 460454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 495834 -7654 496454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 531834 -7654 532454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 567834 -7654 568454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 41514 -7654 42134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 77514 354900 78134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 113514 -7654 114134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 149514 -7654 150134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 185514 354900 186134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 221514 -7654 222134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 257514 27193 258134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 293514 -7654 294134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 329514 -7654 330134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 365514 -7654 366134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 401514 -7654 402134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 437514 -7654 438134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 473514 -7654 474134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 509514 -7654 510134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 545514 -7654 546134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 12954 -7654 13574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 48954 -7654 49574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 84954 -7654 85574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 120954 -7654 121574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 156954 -7654 157574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 192954 -7654 193574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 228954 -7654 229574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 264954 -7654 265574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 300954 -7654 301574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 336954 -7654 337574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 372954 -7654 373574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 408954 -7654 409574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 444954 -7654 445574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 480954 -7654 481574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 516954 -7654 517574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 552954 -7654 553574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal2 s 542 -960 654 480 0 FreeSans 560 90 0 0 wb_clk_i
port 540 nsew
flabel metal2 s 1646 -960 1758 480 0 FreeSans 560 90 0 0 wb_rst_i
port 541 nsew
flabel metal2 s 2842 -960 2954 480 0 FreeSans 560 90 0 0 wbs_ack_o
port 542 nsew
flabel metal2 s 7626 -960 7738 480 0 FreeSans 560 90 0 0 wbs_adr_i[0]
port 543 nsew
flabel metal2 s 47830 -960 47942 480 0 FreeSans 560 90 0 0 wbs_adr_i[10]
port 544 nsew
flabel metal2 s 51326 -960 51438 480 0 FreeSans 560 90 0 0 wbs_adr_i[11]
port 545 nsew
flabel metal2 s 54914 -960 55026 480 0 FreeSans 560 90 0 0 wbs_adr_i[12]
port 546 nsew
flabel metal2 s 58410 -960 58522 480 0 FreeSans 560 90 0 0 wbs_adr_i[13]
port 547 nsew
flabel metal2 s 61998 -960 62110 480 0 FreeSans 560 90 0 0 wbs_adr_i[14]
port 548 nsew
flabel metal2 s 65494 -960 65606 480 0 FreeSans 560 90 0 0 wbs_adr_i[15]
port 549 nsew
flabel metal2 s 69082 -960 69194 480 0 FreeSans 560 90 0 0 wbs_adr_i[16]
port 550 nsew
flabel metal2 s 72578 -960 72690 480 0 FreeSans 560 90 0 0 wbs_adr_i[17]
port 551 nsew
flabel metal2 s 76166 -960 76278 480 0 FreeSans 560 90 0 0 wbs_adr_i[18]
port 552 nsew
flabel metal2 s 79662 -960 79774 480 0 FreeSans 560 90 0 0 wbs_adr_i[19]
port 553 nsew
flabel metal2 s 12318 -960 12430 480 0 FreeSans 560 90 0 0 wbs_adr_i[1]
port 554 nsew
flabel metal2 s 83250 -960 83362 480 0 FreeSans 560 90 0 0 wbs_adr_i[20]
port 555 nsew
flabel metal2 s 86838 -960 86950 480 0 FreeSans 560 90 0 0 wbs_adr_i[21]
port 556 nsew
flabel metal2 s 90334 -960 90446 480 0 FreeSans 560 90 0 0 wbs_adr_i[22]
port 557 nsew
flabel metal2 s 93922 -960 94034 480 0 FreeSans 560 90 0 0 wbs_adr_i[23]
port 558 nsew
flabel metal2 s 97418 -960 97530 480 0 FreeSans 560 90 0 0 wbs_adr_i[24]
port 559 nsew
flabel metal2 s 101006 -960 101118 480 0 FreeSans 560 90 0 0 wbs_adr_i[25]
port 560 nsew
flabel metal2 s 104502 -960 104614 480 0 FreeSans 560 90 0 0 wbs_adr_i[26]
port 561 nsew
flabel metal2 s 108090 -960 108202 480 0 FreeSans 560 90 0 0 wbs_adr_i[27]
port 562 nsew
flabel metal2 s 111586 -960 111698 480 0 FreeSans 560 90 0 0 wbs_adr_i[28]
port 563 nsew
flabel metal2 s 115174 -960 115286 480 0 FreeSans 560 90 0 0 wbs_adr_i[29]
port 564 nsew
flabel metal2 s 17010 -960 17122 480 0 FreeSans 560 90 0 0 wbs_adr_i[2]
port 565 nsew
flabel metal2 s 118762 -960 118874 480 0 FreeSans 560 90 0 0 wbs_adr_i[30]
port 566 nsew
flabel metal2 s 122258 -960 122370 480 0 FreeSans 560 90 0 0 wbs_adr_i[31]
port 567 nsew
flabel metal2 s 21794 -960 21906 480 0 FreeSans 560 90 0 0 wbs_adr_i[3]
port 568 nsew
flabel metal2 s 26486 -960 26598 480 0 FreeSans 560 90 0 0 wbs_adr_i[4]
port 569 nsew
flabel metal2 s 30074 -960 30186 480 0 FreeSans 560 90 0 0 wbs_adr_i[5]
port 570 nsew
flabel metal2 s 33570 -960 33682 480 0 FreeSans 560 90 0 0 wbs_adr_i[6]
port 571 nsew
flabel metal2 s 37158 -960 37270 480 0 FreeSans 560 90 0 0 wbs_adr_i[7]
port 572 nsew
flabel metal2 s 40654 -960 40766 480 0 FreeSans 560 90 0 0 wbs_adr_i[8]
port 573 nsew
flabel metal2 s 44242 -960 44354 480 0 FreeSans 560 90 0 0 wbs_adr_i[9]
port 574 nsew
flabel metal2 s 4038 -960 4150 480 0 FreeSans 560 90 0 0 wbs_cyc_i
port 575 nsew
flabel metal2 s 8730 -960 8842 480 0 FreeSans 560 90 0 0 wbs_dat_i[0]
port 576 nsew
flabel metal2 s 48934 -960 49046 480 0 FreeSans 560 90 0 0 wbs_dat_i[10]
port 577 nsew
flabel metal2 s 52522 -960 52634 480 0 FreeSans 560 90 0 0 wbs_dat_i[11]
port 578 nsew
flabel metal2 s 56018 -960 56130 480 0 FreeSans 560 90 0 0 wbs_dat_i[12]
port 579 nsew
flabel metal2 s 59606 -960 59718 480 0 FreeSans 560 90 0 0 wbs_dat_i[13]
port 580 nsew
flabel metal2 s 63194 -960 63306 480 0 FreeSans 560 90 0 0 wbs_dat_i[14]
port 581 nsew
flabel metal2 s 66690 -960 66802 480 0 FreeSans 560 90 0 0 wbs_dat_i[15]
port 582 nsew
flabel metal2 s 70278 -960 70390 480 0 FreeSans 560 90 0 0 wbs_dat_i[16]
port 583 nsew
flabel metal2 s 73774 -960 73886 480 0 FreeSans 560 90 0 0 wbs_dat_i[17]
port 584 nsew
flabel metal2 s 77362 -960 77474 480 0 FreeSans 560 90 0 0 wbs_dat_i[18]
port 585 nsew
flabel metal2 s 80858 -960 80970 480 0 FreeSans 560 90 0 0 wbs_dat_i[19]
port 586 nsew
flabel metal2 s 13514 -960 13626 480 0 FreeSans 560 90 0 0 wbs_dat_i[1]
port 587 nsew
flabel metal2 s 84446 -960 84558 480 0 FreeSans 560 90 0 0 wbs_dat_i[20]
port 588 nsew
flabel metal2 s 87942 -960 88054 480 0 FreeSans 560 90 0 0 wbs_dat_i[21]
port 589 nsew
flabel metal2 s 91530 -960 91642 480 0 FreeSans 560 90 0 0 wbs_dat_i[22]
port 590 nsew
flabel metal2 s 95118 -960 95230 480 0 FreeSans 560 90 0 0 wbs_dat_i[23]
port 591 nsew
flabel metal2 s 98614 -960 98726 480 0 FreeSans 560 90 0 0 wbs_dat_i[24]
port 592 nsew
flabel metal2 s 102202 -960 102314 480 0 FreeSans 560 90 0 0 wbs_dat_i[25]
port 593 nsew
flabel metal2 s 105698 -960 105810 480 0 FreeSans 560 90 0 0 wbs_dat_i[26]
port 594 nsew
flabel metal2 s 109286 -960 109398 480 0 FreeSans 560 90 0 0 wbs_dat_i[27]
port 595 nsew
flabel metal2 s 112782 -960 112894 480 0 FreeSans 560 90 0 0 wbs_dat_i[28]
port 596 nsew
flabel metal2 s 116370 -960 116482 480 0 FreeSans 560 90 0 0 wbs_dat_i[29]
port 597 nsew
flabel metal2 s 18206 -960 18318 480 0 FreeSans 560 90 0 0 wbs_dat_i[2]
port 598 nsew
flabel metal2 s 119866 -960 119978 480 0 FreeSans 560 90 0 0 wbs_dat_i[30]
port 599 nsew
flabel metal2 s 123454 -960 123566 480 0 FreeSans 560 90 0 0 wbs_dat_i[31]
port 600 nsew
flabel metal2 s 22990 -960 23102 480 0 FreeSans 560 90 0 0 wbs_dat_i[3]
port 601 nsew
flabel metal2 s 27682 -960 27794 480 0 FreeSans 560 90 0 0 wbs_dat_i[4]
port 602 nsew
flabel metal2 s 31270 -960 31382 480 0 FreeSans 560 90 0 0 wbs_dat_i[5]
port 603 nsew
flabel metal2 s 34766 -960 34878 480 0 FreeSans 560 90 0 0 wbs_dat_i[6]
port 604 nsew
flabel metal2 s 38354 -960 38466 480 0 FreeSans 560 90 0 0 wbs_dat_i[7]
port 605 nsew
flabel metal2 s 41850 -960 41962 480 0 FreeSans 560 90 0 0 wbs_dat_i[8]
port 606 nsew
flabel metal2 s 45438 -960 45550 480 0 FreeSans 560 90 0 0 wbs_dat_i[9]
port 607 nsew
flabel metal2 s 9926 -960 10038 480 0 FreeSans 560 90 0 0 wbs_dat_o[0]
port 608 nsew
flabel metal2 s 50130 -960 50242 480 0 FreeSans 560 90 0 0 wbs_dat_o[10]
port 609 nsew
flabel metal2 s 53718 -960 53830 480 0 FreeSans 560 90 0 0 wbs_dat_o[11]
port 610 nsew
flabel metal2 s 57214 -960 57326 480 0 FreeSans 560 90 0 0 wbs_dat_o[12]
port 611 nsew
flabel metal2 s 60802 -960 60914 480 0 FreeSans 560 90 0 0 wbs_dat_o[13]
port 612 nsew
flabel metal2 s 64298 -960 64410 480 0 FreeSans 560 90 0 0 wbs_dat_o[14]
port 613 nsew
flabel metal2 s 67886 -960 67998 480 0 FreeSans 560 90 0 0 wbs_dat_o[15]
port 614 nsew
flabel metal2 s 71474 -960 71586 480 0 FreeSans 560 90 0 0 wbs_dat_o[16]
port 615 nsew
flabel metal2 s 74970 -960 75082 480 0 FreeSans 560 90 0 0 wbs_dat_o[17]
port 616 nsew
flabel metal2 s 78558 -960 78670 480 0 FreeSans 560 90 0 0 wbs_dat_o[18]
port 617 nsew
flabel metal2 s 82054 -960 82166 480 0 FreeSans 560 90 0 0 wbs_dat_o[19]
port 618 nsew
flabel metal2 s 14710 -960 14822 480 0 FreeSans 560 90 0 0 wbs_dat_o[1]
port 619 nsew
flabel metal2 s 85642 -960 85754 480 0 FreeSans 560 90 0 0 wbs_dat_o[20]
port 620 nsew
flabel metal2 s 89138 -960 89250 480 0 FreeSans 560 90 0 0 wbs_dat_o[21]
port 621 nsew
flabel metal2 s 92726 -960 92838 480 0 FreeSans 560 90 0 0 wbs_dat_o[22]
port 622 nsew
flabel metal2 s 96222 -960 96334 480 0 FreeSans 560 90 0 0 wbs_dat_o[23]
port 623 nsew
flabel metal2 s 99810 -960 99922 480 0 FreeSans 560 90 0 0 wbs_dat_o[24]
port 624 nsew
flabel metal2 s 103306 -960 103418 480 0 FreeSans 560 90 0 0 wbs_dat_o[25]
port 625 nsew
flabel metal2 s 106894 -960 107006 480 0 FreeSans 560 90 0 0 wbs_dat_o[26]
port 626 nsew
flabel metal2 s 110482 -960 110594 480 0 FreeSans 560 90 0 0 wbs_dat_o[27]
port 627 nsew
flabel metal2 s 113978 -960 114090 480 0 FreeSans 560 90 0 0 wbs_dat_o[28]
port 628 nsew
flabel metal2 s 117566 -960 117678 480 0 FreeSans 560 90 0 0 wbs_dat_o[29]
port 629 nsew
flabel metal2 s 19402 -960 19514 480 0 FreeSans 560 90 0 0 wbs_dat_o[2]
port 630 nsew
flabel metal2 s 121062 -960 121174 480 0 FreeSans 560 90 0 0 wbs_dat_o[30]
port 631 nsew
flabel metal2 s 124650 -960 124762 480 0 FreeSans 560 90 0 0 wbs_dat_o[31]
port 632 nsew
flabel metal2 s 24186 -960 24298 480 0 FreeSans 560 90 0 0 wbs_dat_o[3]
port 633 nsew
flabel metal2 s 28878 -960 28990 480 0 FreeSans 560 90 0 0 wbs_dat_o[4]
port 634 nsew
flabel metal2 s 32374 -960 32486 480 0 FreeSans 560 90 0 0 wbs_dat_o[5]
port 635 nsew
flabel metal2 s 35962 -960 36074 480 0 FreeSans 560 90 0 0 wbs_dat_o[6]
port 636 nsew
flabel metal2 s 39550 -960 39662 480 0 FreeSans 560 90 0 0 wbs_dat_o[7]
port 637 nsew
flabel metal2 s 43046 -960 43158 480 0 FreeSans 560 90 0 0 wbs_dat_o[8]
port 638 nsew
flabel metal2 s 46634 -960 46746 480 0 FreeSans 560 90 0 0 wbs_dat_o[9]
port 639 nsew
flabel metal2 s 11122 -960 11234 480 0 FreeSans 560 90 0 0 wbs_sel_i[0]
port 640 nsew
flabel metal2 s 15906 -960 16018 480 0 FreeSans 560 90 0 0 wbs_sel_i[1]
port 641 nsew
flabel metal2 s 20598 -960 20710 480 0 FreeSans 560 90 0 0 wbs_sel_i[2]
port 642 nsew
flabel metal2 s 25290 -960 25402 480 0 FreeSans 560 90 0 0 wbs_sel_i[3]
port 643 nsew
flabel metal2 s 5234 -960 5346 480 0 FreeSans 560 90 0 0 wbs_stb_i
port 644 nsew
flabel metal2 s 6430 -960 6542 480 0 FreeSans 560 90 0 0 wbs_we_i
port 645 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
